module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg,
    VDD,
    VSS);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;
 inout VDD;
 inout VSS;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire _482_;
 wire _483_;
 wire _484_;
 wire _485_;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;

 INV_X1 _486_ (.A(\dpath.a_lt_b$in1[11] ),
    .ZN(_036_));
 INV_X1 _487_ (.A(\dpath.a_lt_b$in1[10] ),
    .ZN(_037_));
 INV_X2 _488_ (.A(\dpath.a_lt_b$in1[9] ),
    .ZN(_038_));
 INV_X2 _489_ (.A(\dpath.a_lt_b$in1[8] ),
    .ZN(_039_));
 NAND4_X1 _490_ (.A1(_036_),
    .A2(_037_),
    .A3(_038_),
    .A4(_039_),
    .ZN(_040_));
 INV_X1 _491_ (.A(\dpath.a_lt_b$in1[15] ),
    .ZN(_041_));
 INV_X2 _492_ (.A(\dpath.a_lt_b$in1[14] ),
    .ZN(_042_));
 INV_X1 _493_ (.A(\dpath.a_lt_b$in1[13] ),
    .ZN(_043_));
 INV_X2 _494_ (.A(\dpath.a_lt_b$in1[12] ),
    .ZN(_044_));
 NAND4_X1 _495_ (.A1(_041_),
    .A2(_042_),
    .A3(_043_),
    .A4(_044_),
    .ZN(_045_));
 INV_X2 _496_ (.A(\dpath.a_lt_b$in1[3] ),
    .ZN(_046_));
 INV_X2 _497_ (.A(\dpath.a_lt_b$in1[2] ),
    .ZN(_047_));
 INV_X2 _498_ (.A(\dpath.a_lt_b$in1[1] ),
    .ZN(_048_));
 INV_X2 _499_ (.A(\dpath.a_lt_b$in1[0] ),
    .ZN(_049_));
 NAND4_X1 _500_ (.A1(_046_),
    .A2(_047_),
    .A3(_048_),
    .A4(_049_),
    .ZN(_050_));
 INV_X2 _501_ (.A(\dpath.a_lt_b$in1[7] ),
    .ZN(_051_));
 INV_X2 _502_ (.A(\dpath.a_lt_b$in1[6] ),
    .ZN(_052_));
 INV_X2 _503_ (.A(\dpath.a_lt_b$in1[5] ),
    .ZN(_053_));
 INV_X1 _504_ (.A(\dpath.a_lt_b$in1[4] ),
    .ZN(_054_));
 NAND4_X1 _505_ (.A1(_051_),
    .A2(_052_),
    .A3(_053_),
    .A4(_054_),
    .ZN(_055_));
 NOR4_X1 _506_ (.A1(_040_),
    .A2(_045_),
    .A3(_050_),
    .A4(_055_),
    .ZN(_056_));
 BUF_X1 _507_ (.A(\ctrl.state.out[2] ),
    .Z(_057_));
 INV_X1 _508_ (.A(_057_),
    .ZN(_058_));
 OR2_X1 _509_ (.A1(_058_),
    .A2(reset),
    .ZN(_059_));
 BUF_X1 _510_ (.A(req_rdy),
    .Z(_060_));
 BUF_X1 _511_ (.A(_060_),
    .Z(_061_));
 BUF_X1 _512_ (.A(_061_),
    .Z(_062_));
 NAND2_X1 _513_ (.A1(_062_),
    .A2(req_val),
    .ZN(_063_));
 OAI22_X1 _514_ (.A1(_056_),
    .A2(_059_),
    .B1(reset),
    .B2(_063_),
    .ZN(_002_));
 BUF_X2 _515_ (.A(_003_),
    .Z(_064_));
 AND3_X1 _516_ (.A1(_058_),
    .A2(\ctrl.state.out[1] ),
    .A3(_064_),
    .ZN(resp_val));
 AOI21_X1 _517_ (.A(reset),
    .B1(resp_val),
    .B2(resp_rdy),
    .ZN(_065_));
 BUF_X1 _518_ (.A(_060_),
    .Z(_066_));
 BUF_X1 _519_ (.A(_066_),
    .Z(_067_));
 INV_X1 _520_ (.A(_067_),
    .ZN(_068_));
 OAI21_X1 _521_ (.A(_065_),
    .B1(_068_),
    .B2(req_val),
    .ZN(_000_));
 NAND2_X1 _522_ (.A1(_065_),
    .A2(\ctrl.state.out[1] ),
    .ZN(_069_));
 INV_X1 _523_ (.A(_056_),
    .ZN(_070_));
 OAI21_X1 _524_ (.A(_069_),
    .B1(_070_),
    .B2(_059_),
    .ZN(_001_));
 XNOR2_X1 _525_ (.A(_049_),
    .B(\dpath.a_lt_b$in0[0] ),
    .ZN(resp_msg[0]));
 BUF_X2 _526_ (.A(\dpath.a_lt_b$in0[1] ),
    .Z(_071_));
 NAND2_X1 _527_ (.A1(_048_),
    .A2(_071_),
    .ZN(_072_));
 NOR2_X1 _528_ (.A1(_049_),
    .A2(\dpath.a_lt_b$in0[0] ),
    .ZN(_073_));
 NOR2_X1 _529_ (.A1(_048_),
    .A2(_071_),
    .ZN(_074_));
 OAI21_X1 _530_ (.A(_072_),
    .B1(_073_),
    .B2(_074_),
    .ZN(_075_));
 NAND2_X1 _531_ (.A1(_046_),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_076_));
 INV_X1 _532_ (.A(\dpath.a_lt_b$in0[3] ),
    .ZN(_077_));
 NAND2_X1 _533_ (.A1(_077_),
    .A2(\dpath.a_lt_b$in1[3] ),
    .ZN(_078_));
 NAND2_X2 _534_ (.A1(_076_),
    .A2(_078_),
    .ZN(_079_));
 NAND2_X1 _535_ (.A1(_047_),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_080_));
 INV_X1 _536_ (.A(\dpath.a_lt_b$in0[2] ),
    .ZN(_081_));
 NAND2_X1 _537_ (.A1(_081_),
    .A2(\dpath.a_lt_b$in1[2] ),
    .ZN(_082_));
 NAND2_X2 _538_ (.A1(_080_),
    .A2(_082_),
    .ZN(_083_));
 NOR2_X2 _539_ (.A1(_079_),
    .A2(_083_),
    .ZN(_084_));
 NAND2_X1 _540_ (.A1(_075_),
    .A2(_084_),
    .ZN(_085_));
 NOR2_X1 _541_ (.A1(_046_),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_086_));
 OAI21_X1 _542_ (.A(_076_),
    .B1(_086_),
    .B2(_080_),
    .ZN(_087_));
 INV_X1 _543_ (.A(_087_),
    .ZN(_088_));
 NAND2_X2 _544_ (.A1(_085_),
    .A2(_088_),
    .ZN(_089_));
 INV_X1 _545_ (.A(\dpath.a_lt_b$in0[7] ),
    .ZN(_090_));
 NAND2_X2 _546_ (.A1(_090_),
    .A2(\dpath.a_lt_b$in1[7] ),
    .ZN(_091_));
 NAND2_X2 _547_ (.A1(_051_),
    .A2(\dpath.a_lt_b$in0[7] ),
    .ZN(_092_));
 NAND2_X2 _548_ (.A1(_091_),
    .A2(_092_),
    .ZN(_093_));
 NAND2_X2 _549_ (.A1(_052_),
    .A2(\dpath.a_lt_b$in0[6] ),
    .ZN(_094_));
 INV_X1 _550_ (.A(\dpath.a_lt_b$in0[6] ),
    .ZN(_095_));
 NAND2_X2 _551_ (.A1(_095_),
    .A2(\dpath.a_lt_b$in1[6] ),
    .ZN(_096_));
 NAND2_X4 _552_ (.A1(_094_),
    .A2(_096_),
    .ZN(_097_));
 NOR2_X4 _553_ (.A1(_093_),
    .A2(_097_),
    .ZN(_098_));
 NAND2_X2 _554_ (.A1(_053_),
    .A2(\dpath.a_lt_b$in0[5] ),
    .ZN(_099_));
 INV_X1 _555_ (.A(\dpath.a_lt_b$in0[5] ),
    .ZN(_100_));
 NAND2_X2 _556_ (.A1(_100_),
    .A2(\dpath.a_lt_b$in1[5] ),
    .ZN(_101_));
 NAND2_X2 _557_ (.A1(_099_),
    .A2(_101_),
    .ZN(_102_));
 NAND2_X1 _558_ (.A1(_054_),
    .A2(\dpath.a_lt_b$in0[4] ),
    .ZN(_103_));
 INV_X1 _559_ (.A(\dpath.a_lt_b$in0[4] ),
    .ZN(_104_));
 NAND2_X1 _560_ (.A1(_104_),
    .A2(\dpath.a_lt_b$in1[4] ),
    .ZN(_105_));
 NAND2_X2 _561_ (.A1(_103_),
    .A2(_105_),
    .ZN(_106_));
 NOR2_X2 _562_ (.A1(_102_),
    .A2(_106_),
    .ZN(_107_));
 AND2_X2 _563_ (.A1(_098_),
    .A2(_107_),
    .ZN(_108_));
 NAND2_X2 _564_ (.A1(_089_),
    .A2(_108_),
    .ZN(_109_));
 NAND2_X1 _565_ (.A1(_092_),
    .A2(_094_),
    .ZN(_110_));
 NAND2_X2 _566_ (.A1(_110_),
    .A2(_091_),
    .ZN(_111_));
 INV_X1 _567_ (.A(_111_),
    .ZN(_112_));
 INV_X1 _568_ (.A(_099_),
    .ZN(_113_));
 NOR2_X1 _569_ (.A1(_104_),
    .A2(\dpath.a_lt_b$in1[4] ),
    .ZN(_114_));
 OAI21_X2 _570_ (.A(_101_),
    .B1(_113_),
    .B2(_114_),
    .ZN(_115_));
 INV_X1 _571_ (.A(_115_),
    .ZN(_116_));
 AOI21_X4 _572_ (.A(_112_),
    .B1(_116_),
    .B2(_098_),
    .ZN(_117_));
 NAND2_X4 _573_ (.A1(_109_),
    .A2(_117_),
    .ZN(_118_));
 INV_X1 _574_ (.A(\dpath.a_lt_b$in0[13] ),
    .ZN(_119_));
 NOR2_X2 _575_ (.A1(_119_),
    .A2(\dpath.a_lt_b$in1[13] ),
    .ZN(_120_));
 INV_X1 _576_ (.A(_120_),
    .ZN(_121_));
 NAND2_X1 _577_ (.A1(_119_),
    .A2(\dpath.a_lt_b$in1[13] ),
    .ZN(_122_));
 NAND2_X2 _578_ (.A1(_121_),
    .A2(_122_),
    .ZN(_123_));
 INV_X2 _579_ (.A(_123_),
    .ZN(_124_));
 INV_X1 _580_ (.A(\dpath.a_lt_b$in0[12] ),
    .ZN(_125_));
 NOR2_X2 _581_ (.A1(_125_),
    .A2(\dpath.a_lt_b$in1[12] ),
    .ZN(_126_));
 NOR2_X2 _582_ (.A1(_044_),
    .A2(\dpath.a_lt_b$in0[12] ),
    .ZN(_127_));
 NOR2_X4 _583_ (.A1(_126_),
    .A2(_127_),
    .ZN(_128_));
 NAND2_X1 _584_ (.A1(_124_),
    .A2(_128_),
    .ZN(_129_));
 NAND2_X2 _585_ (.A1(_042_),
    .A2(\dpath.a_lt_b$in0[14] ),
    .ZN(_130_));
 INV_X1 _586_ (.A(\dpath.a_lt_b$in0[14] ),
    .ZN(_131_));
 NAND2_X1 _587_ (.A1(_131_),
    .A2(\dpath.a_lt_b$in1[14] ),
    .ZN(_132_));
 NAND2_X2 _588_ (.A1(_130_),
    .A2(_132_),
    .ZN(_133_));
 INV_X2 _589_ (.A(_133_),
    .ZN(_134_));
 XNOR2_X1 _590_ (.A(\dpath.a_lt_b$in1[15] ),
    .B(\dpath.a_lt_b$in0[15] ),
    .ZN(_135_));
 NAND2_X1 _591_ (.A1(_134_),
    .A2(_135_),
    .ZN(_136_));
 NOR2_X2 _592_ (.A1(_129_),
    .A2(_136_),
    .ZN(_137_));
 NAND2_X1 _593_ (.A1(_036_),
    .A2(\dpath.a_lt_b$in0[11] ),
    .ZN(_138_));
 INV_X1 _594_ (.A(\dpath.a_lt_b$in0[11] ),
    .ZN(_139_));
 NAND2_X1 _595_ (.A1(_139_),
    .A2(\dpath.a_lt_b$in1[11] ),
    .ZN(_140_));
 NAND2_X2 _596_ (.A1(_138_),
    .A2(_140_),
    .ZN(_141_));
 NAND2_X2 _597_ (.A1(_037_),
    .A2(\dpath.a_lt_b$in0[10] ),
    .ZN(_142_));
 INV_X1 _598_ (.A(\dpath.a_lt_b$in0[10] ),
    .ZN(_143_));
 NAND2_X1 _599_ (.A1(_143_),
    .A2(\dpath.a_lt_b$in1[10] ),
    .ZN(_144_));
 NAND2_X2 _600_ (.A1(_142_),
    .A2(_144_),
    .ZN(_145_));
 NOR2_X4 _601_ (.A1(_141_),
    .A2(_145_),
    .ZN(_146_));
 INV_X1 _602_ (.A(_146_),
    .ZN(_147_));
 NAND2_X4 _603_ (.A1(_038_),
    .A2(\dpath.a_lt_b$in0[9] ),
    .ZN(_148_));
 INV_X1 _604_ (.A(\dpath.a_lt_b$in0[9] ),
    .ZN(_149_));
 NAND2_X2 _605_ (.A1(_149_),
    .A2(\dpath.a_lt_b$in1[9] ),
    .ZN(_150_));
 NAND2_X2 _606_ (.A1(_148_),
    .A2(_150_),
    .ZN(_151_));
 INV_X2 _607_ (.A(_151_),
    .ZN(_152_));
 NAND2_X2 _608_ (.A1(_039_),
    .A2(\dpath.a_lt_b$in0[8] ),
    .ZN(_153_));
 INV_X1 _609_ (.A(\dpath.a_lt_b$in0[8] ),
    .ZN(_154_));
 NAND2_X1 _610_ (.A1(_154_),
    .A2(\dpath.a_lt_b$in1[8] ),
    .ZN(_155_));
 NAND2_X2 _611_ (.A1(_153_),
    .A2(_155_),
    .ZN(_156_));
 INV_X4 _612_ (.A(_156_),
    .ZN(_157_));
 NAND2_X2 _613_ (.A1(_152_),
    .A2(_157_),
    .ZN(_158_));
 NOR2_X2 _614_ (.A1(_147_),
    .A2(_158_),
    .ZN(_159_));
 AND2_X2 _615_ (.A1(_137_),
    .A2(_159_),
    .ZN(_160_));
 NAND2_X4 _616_ (.A1(_118_),
    .A2(_160_),
    .ZN(_161_));
 NAND2_X1 _617_ (.A1(_148_),
    .A2(_153_),
    .ZN(_162_));
 NAND2_X1 _618_ (.A1(_162_),
    .A2(_150_),
    .ZN(_163_));
 INV_X1 _619_ (.A(_163_),
    .ZN(_164_));
 NAND2_X2 _620_ (.A1(_146_),
    .A2(_164_),
    .ZN(_165_));
 INV_X1 _621_ (.A(_138_),
    .ZN(_166_));
 INV_X1 _622_ (.A(_142_),
    .ZN(_167_));
 OAI21_X1 _623_ (.A(_140_),
    .B1(_166_),
    .B2(_167_),
    .ZN(_168_));
 NAND2_X1 _624_ (.A1(_165_),
    .A2(_168_),
    .ZN(_169_));
 NAND2_X1 _625_ (.A1(_169_),
    .A2(_137_),
    .ZN(_170_));
 OAI21_X1 _626_ (.A(_122_),
    .B1(_120_),
    .B2(_126_),
    .ZN(_171_));
 NOR2_X1 _627_ (.A1(_171_),
    .A2(_136_),
    .ZN(_172_));
 NAND2_X1 _628_ (.A1(_041_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .ZN(_173_));
 INV_X1 _629_ (.A(_135_),
    .ZN(_174_));
 OAI21_X1 _630_ (.A(_173_),
    .B1(_174_),
    .B2(_130_),
    .ZN(_175_));
 NOR2_X1 _631_ (.A1(_172_),
    .A2(_175_),
    .ZN(_176_));
 NAND2_X1 _632_ (.A1(_170_),
    .A2(_176_),
    .ZN(_177_));
 INV_X4 _633_ (.A(_177_),
    .ZN(_178_));
 NAND2_X4 _634_ (.A1(_161_),
    .A2(_178_),
    .ZN(_179_));
 NAND2_X1 _635_ (.A1(_057_),
    .A2(_003_),
    .ZN(_180_));
 INV_X1 _636_ (.A(_180_),
    .ZN(_181_));
 NAND3_X1 _637_ (.A1(_179_),
    .A2(resp_msg[0]),
    .A3(_181_),
    .ZN(_182_));
 NAND4_X4 _638_ (.A1(_161_),
    .A2(_057_),
    .A3(_064_),
    .A4(_178_),
    .ZN(_183_));
 OAI21_X1 _639_ (.A(_182_),
    .B1(_183_),
    .B2(_049_),
    .ZN(_184_));
 NOR2_X1 _640_ (.A1(_058_),
    .A2(_060_),
    .ZN(_185_));
 BUF_X2 _641_ (.A(_185_),
    .Z(_186_));
 NAND2_X1 _642_ (.A1(_184_),
    .A2(_186_),
    .ZN(_187_));
 NOR2_X1 _643_ (.A1(_060_),
    .A2(_057_),
    .ZN(_188_));
 BUF_X1 _644_ (.A(_188_),
    .Z(_189_));
 AND2_X1 _645_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[0] ),
    .ZN(_190_));
 AOI21_X1 _646_ (.A(_190_),
    .B1(_067_),
    .B2(req_msg[16]),
    .ZN(_191_));
 NAND2_X1 _647_ (.A1(_187_),
    .A2(_191_),
    .ZN(_004_));
 NAND3_X4 _648_ (.A1(_161_),
    .A2(_057_),
    .A3(_178_),
    .ZN(_192_));
 INV_X2 _649_ (.A(_192_),
    .ZN(_193_));
 NAND3_X1 _650_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[10] ),
    .A3(_064_),
    .ZN(_194_));
 NAND2_X1 _651_ (.A1(_107_),
    .A2(_087_),
    .ZN(_195_));
 NAND2_X1 _652_ (.A1(_195_),
    .A2(_115_),
    .ZN(_196_));
 INV_X1 _653_ (.A(_196_),
    .ZN(_197_));
 NAND3_X1 _654_ (.A1(_075_),
    .A2(_084_),
    .A3(_107_),
    .ZN(_198_));
 NAND2_X2 _655_ (.A1(_197_),
    .A2(_198_),
    .ZN(_199_));
 NAND3_X1 _656_ (.A1(_098_),
    .A2(_152_),
    .A3(_157_),
    .ZN(_200_));
 INV_X1 _657_ (.A(_200_),
    .ZN(_201_));
 NAND2_X1 _658_ (.A1(_199_),
    .A2(_201_),
    .ZN(_202_));
 OAI21_X1 _659_ (.A(_163_),
    .B1(_158_),
    .B2(_111_),
    .ZN(_203_));
 INV_X1 _660_ (.A(_203_),
    .ZN(_204_));
 NAND2_X1 _661_ (.A1(_202_),
    .A2(_204_),
    .ZN(_205_));
 XNOR2_X1 _662_ (.A(_205_),
    .B(_145_),
    .ZN(resp_msg[10]));
 AOI21_X4 _663_ (.A(_180_),
    .B1(_161_),
    .B2(_178_),
    .ZN(_206_));
 NAND2_X1 _664_ (.A1(resp_msg[10]),
    .A2(_206_),
    .ZN(_207_));
 NAND2_X1 _665_ (.A1(_194_),
    .A2(_207_),
    .ZN(_208_));
 NAND2_X1 _666_ (.A1(_208_),
    .A2(_186_),
    .ZN(_209_));
 AND2_X1 _667_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[10] ),
    .ZN(_210_));
 AOI21_X1 _668_ (.A(_210_),
    .B1(_067_),
    .B2(req_msg[26]),
    .ZN(_211_));
 NAND2_X1 _669_ (.A1(_209_),
    .A2(_211_),
    .ZN(_005_));
 NAND3_X1 _670_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[11] ),
    .A3(_064_),
    .ZN(_212_));
 INV_X1 _671_ (.A(_083_),
    .ZN(_213_));
 XNOR2_X1 _672_ (.A(\dpath.a_lt_b$in1[1] ),
    .B(_071_),
    .ZN(_214_));
 INV_X1 _673_ (.A(_073_),
    .ZN(_215_));
 NAND3_X1 _674_ (.A1(_213_),
    .A2(_214_),
    .A3(_215_),
    .ZN(_216_));
 NOR2_X1 _675_ (.A1(_047_),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_217_));
 OAI21_X1 _676_ (.A(_080_),
    .B1(_217_),
    .B2(_072_),
    .ZN(_218_));
 INV_X1 _677_ (.A(_218_),
    .ZN(_219_));
 NAND2_X2 _678_ (.A1(_216_),
    .A2(_219_),
    .ZN(_220_));
 NOR2_X2 _679_ (.A1(_079_),
    .A2(_106_),
    .ZN(_221_));
 INV_X1 _680_ (.A(_221_),
    .ZN(_222_));
 NOR2_X4 _681_ (.A1(_097_),
    .A2(_102_),
    .ZN(_223_));
 INV_X1 _682_ (.A(_223_),
    .ZN(_224_));
 NOR2_X2 _683_ (.A1(_222_),
    .A2(_224_),
    .ZN(_225_));
 NAND2_X2 _684_ (.A1(_220_),
    .A2(_225_),
    .ZN(_226_));
 NAND2_X1 _685_ (.A1(_094_),
    .A2(_099_),
    .ZN(_227_));
 NAND2_X1 _686_ (.A1(_227_),
    .A2(_096_),
    .ZN(_228_));
 INV_X1 _687_ (.A(_228_),
    .ZN(_229_));
 INV_X1 _688_ (.A(_076_),
    .ZN(_230_));
 OAI21_X2 _689_ (.A(_105_),
    .B1(_230_),
    .B2(_114_),
    .ZN(_231_));
 INV_X1 _690_ (.A(_231_),
    .ZN(_232_));
 AOI21_X2 _691_ (.A(_229_),
    .B1(_232_),
    .B2(_223_),
    .ZN(_233_));
 NAND2_X4 _692_ (.A1(_226_),
    .A2(_233_),
    .ZN(_234_));
 INV_X1 _693_ (.A(_145_),
    .ZN(_235_));
 NAND2_X2 _694_ (.A1(_235_),
    .A2(_152_),
    .ZN(_236_));
 INV_X1 _695_ (.A(_236_),
    .ZN(_237_));
 INV_X2 _696_ (.A(_093_),
    .ZN(_238_));
 NAND2_X2 _697_ (.A1(_238_),
    .A2(_157_),
    .ZN(_239_));
 INV_X1 _698_ (.A(_239_),
    .ZN(_240_));
 NAND2_X1 _699_ (.A1(_237_),
    .A2(_240_),
    .ZN(_241_));
 INV_X2 _700_ (.A(_241_),
    .ZN(_242_));
 NAND2_X2 _701_ (.A1(_234_),
    .A2(_242_),
    .ZN(_243_));
 INV_X1 _702_ (.A(_148_),
    .ZN(_244_));
 OAI21_X1 _703_ (.A(_144_),
    .B1(_167_),
    .B2(_244_),
    .ZN(_245_));
 NAND2_X1 _704_ (.A1(_092_),
    .A2(_153_),
    .ZN(_246_));
 NAND2_X1 _705_ (.A1(_246_),
    .A2(_155_),
    .ZN(_247_));
 OAI21_X1 _706_ (.A(_245_),
    .B1(_236_),
    .B2(_247_),
    .ZN(_248_));
 INV_X1 _707_ (.A(_248_),
    .ZN(_249_));
 NAND2_X1 _708_ (.A1(_243_),
    .A2(_249_),
    .ZN(_250_));
 NAND2_X1 _709_ (.A1(_250_),
    .A2(_141_),
    .ZN(_251_));
 INV_X1 _710_ (.A(_141_),
    .ZN(_252_));
 NAND3_X1 _711_ (.A1(_243_),
    .A2(_252_),
    .A3(_249_),
    .ZN(_253_));
 NAND2_X1 _712_ (.A1(_251_),
    .A2(_253_),
    .ZN(resp_msg[11]));
 NAND2_X1 _713_ (.A1(resp_msg[11]),
    .A2(_206_),
    .ZN(_254_));
 NAND2_X1 _714_ (.A1(_212_),
    .A2(_254_),
    .ZN(_255_));
 NAND2_X1 _715_ (.A1(_255_),
    .A2(_186_),
    .ZN(_256_));
 AND2_X1 _716_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[11] ),
    .ZN(_257_));
 AOI21_X1 _717_ (.A(_257_),
    .B1(_067_),
    .B2(req_msg[27]),
    .ZN(_258_));
 NAND2_X1 _718_ (.A1(_256_),
    .A2(_258_),
    .ZN(_006_));
 NAND3_X1 _719_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[12] ),
    .A3(_064_),
    .ZN(_259_));
 INV_X1 _720_ (.A(_098_),
    .ZN(_260_));
 OAI21_X1 _721_ (.A(_111_),
    .B1(_260_),
    .B2(_115_),
    .ZN(_261_));
 NAND2_X1 _722_ (.A1(_261_),
    .A2(_159_),
    .ZN(_262_));
 INV_X1 _723_ (.A(_169_),
    .ZN(_263_));
 NAND2_X1 _724_ (.A1(_262_),
    .A2(_263_),
    .ZN(_264_));
 NAND2_X1 _725_ (.A1(_108_),
    .A2(_159_),
    .ZN(_265_));
 INV_X1 _726_ (.A(_089_),
    .ZN(_266_));
 NOR2_X1 _727_ (.A1(_265_),
    .A2(_266_),
    .ZN(_267_));
 NOR2_X1 _728_ (.A1(_264_),
    .A2(_267_),
    .ZN(_268_));
 NAND2_X1 _729_ (.A1(_268_),
    .A2(_128_),
    .ZN(_269_));
 INV_X1 _730_ (.A(_128_),
    .ZN(_270_));
 OAI21_X1 _731_ (.A(_270_),
    .B1(_264_),
    .B2(_267_),
    .ZN(_271_));
 NAND2_X1 _732_ (.A1(_269_),
    .A2(_271_),
    .ZN(resp_msg[12]));
 NAND2_X1 _733_ (.A1(resp_msg[12]),
    .A2(_206_),
    .ZN(_272_));
 NAND2_X1 _734_ (.A1(_259_),
    .A2(_272_),
    .ZN(_273_));
 NAND2_X1 _735_ (.A1(_273_),
    .A2(_186_),
    .ZN(_274_));
 AND2_X1 _736_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[12] ),
    .ZN(_275_));
 AOI21_X1 _737_ (.A(_275_),
    .B1(_067_),
    .B2(req_msg[28]),
    .ZN(_276_));
 NAND2_X1 _738_ (.A1(_274_),
    .A2(_276_),
    .ZN(_007_));
 NAND3_X1 _739_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[13] ),
    .A3(_064_),
    .ZN(_277_));
 NOR2_X2 _740_ (.A1(_270_),
    .A2(_141_),
    .ZN(_278_));
 INV_X1 _741_ (.A(_278_),
    .ZN(_279_));
 NOR2_X2 _742_ (.A1(_279_),
    .A2(_236_),
    .ZN(_280_));
 NOR2_X2 _743_ (.A1(_224_),
    .A2(_239_),
    .ZN(_281_));
 AND2_X1 _744_ (.A1(_280_),
    .A2(_281_),
    .ZN(_282_));
 NAND2_X1 _745_ (.A1(_220_),
    .A2(_221_),
    .ZN(_283_));
 NAND2_X1 _746_ (.A1(_283_),
    .A2(_231_),
    .ZN(_284_));
 NAND2_X1 _747_ (.A1(_282_),
    .A2(_284_),
    .ZN(_285_));
 OAI21_X1 _748_ (.A(_247_),
    .B1(_239_),
    .B2(_228_),
    .ZN(_286_));
 NAND2_X1 _749_ (.A1(_280_),
    .A2(_286_),
    .ZN(_287_));
 INV_X1 _750_ (.A(_127_),
    .ZN(_288_));
 OAI21_X1 _751_ (.A(_288_),
    .B1(_166_),
    .B2(_126_),
    .ZN(_289_));
 INV_X1 _752_ (.A(_289_),
    .ZN(_290_));
 INV_X1 _753_ (.A(_245_),
    .ZN(_291_));
 AOI21_X1 _754_ (.A(_290_),
    .B1(_291_),
    .B2(_278_),
    .ZN(_292_));
 NAND2_X1 _755_ (.A1(_287_),
    .A2(_292_),
    .ZN(_293_));
 INV_X1 _756_ (.A(_293_),
    .ZN(_294_));
 NAND2_X1 _757_ (.A1(_285_),
    .A2(_294_),
    .ZN(_295_));
 NAND2_X1 _758_ (.A1(_295_),
    .A2(_123_),
    .ZN(_296_));
 NAND3_X1 _759_ (.A1(_285_),
    .A2(_294_),
    .A3(_124_),
    .ZN(_297_));
 NAND2_X2 _760_ (.A1(_296_),
    .A2(_297_),
    .ZN(resp_msg[13]));
 NAND2_X1 _761_ (.A1(resp_msg[13]),
    .A2(_206_),
    .ZN(_298_));
 NAND2_X1 _762_ (.A1(_277_),
    .A2(_298_),
    .ZN(_299_));
 NAND2_X1 _763_ (.A1(_299_),
    .A2(_186_),
    .ZN(_300_));
 AND2_X1 _764_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[13] ),
    .ZN(_301_));
 AOI21_X1 _765_ (.A(_301_),
    .B1(_067_),
    .B2(req_msg[29]),
    .ZN(_302_));
 NAND2_X1 _766_ (.A1(_300_),
    .A2(_302_),
    .ZN(_008_));
 NAND3_X1 _767_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[14] ),
    .A3(_064_),
    .ZN(_303_));
 NAND3_X1 _768_ (.A1(_146_),
    .A2(_124_),
    .A3(_128_),
    .ZN(_304_));
 NOR2_X1 _769_ (.A1(_200_),
    .A2(_304_),
    .ZN(_305_));
 NAND2_X1 _770_ (.A1(_199_),
    .A2(_305_),
    .ZN(_306_));
 INV_X1 _771_ (.A(_306_),
    .ZN(_307_));
 INV_X1 _772_ (.A(_304_),
    .ZN(_308_));
 NAND2_X1 _773_ (.A1(_203_),
    .A2(_308_),
    .ZN(_309_));
 NOR2_X1 _774_ (.A1(_129_),
    .A2(_168_),
    .ZN(_310_));
 INV_X1 _775_ (.A(_171_),
    .ZN(_311_));
 NOR2_X1 _776_ (.A1(_310_),
    .A2(_311_),
    .ZN(_312_));
 NAND2_X1 _777_ (.A1(_309_),
    .A2(_312_),
    .ZN(_313_));
 OAI21_X1 _778_ (.A(_133_),
    .B1(_307_),
    .B2(_313_),
    .ZN(_314_));
 INV_X1 _779_ (.A(_313_),
    .ZN(_315_));
 NAND3_X1 _780_ (.A1(_315_),
    .A2(_306_),
    .A3(_134_),
    .ZN(_316_));
 NAND2_X1 _781_ (.A1(_314_),
    .A2(_316_),
    .ZN(resp_msg[14]));
 NAND2_X1 _782_ (.A1(resp_msg[14]),
    .A2(_206_),
    .ZN(_317_));
 NAND2_X1 _783_ (.A1(_303_),
    .A2(_317_),
    .ZN(_318_));
 NAND2_X1 _784_ (.A1(_318_),
    .A2(_186_),
    .ZN(_319_));
 AND2_X1 _785_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[14] ),
    .ZN(_320_));
 AOI21_X1 _786_ (.A(_320_),
    .B1(_067_),
    .B2(req_msg[30]),
    .ZN(_321_));
 NAND2_X1 _787_ (.A1(_319_),
    .A2(_321_),
    .ZN(_009_));
 NAND3_X1 _788_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[15] ),
    .A3(_064_),
    .ZN(_322_));
 NOR2_X1 _789_ (.A1(_123_),
    .A2(_133_),
    .ZN(_323_));
 AND2_X1 _790_ (.A1(_278_),
    .A2(_323_),
    .ZN(_324_));
 AND2_X1 _791_ (.A1(_324_),
    .A2(_242_),
    .ZN(_325_));
 NAND2_X1 _792_ (.A1(_234_),
    .A2(_325_),
    .ZN(_326_));
 NAND2_X1 _793_ (.A1(_324_),
    .A2(_248_),
    .ZN(_327_));
 OAI21_X1 _794_ (.A(_130_),
    .B1(_133_),
    .B2(_121_),
    .ZN(_328_));
 AOI21_X1 _795_ (.A(_328_),
    .B1(_290_),
    .B2(_323_),
    .ZN(_329_));
 NAND2_X1 _796_ (.A1(_327_),
    .A2(_329_),
    .ZN(_330_));
 INV_X1 _797_ (.A(_330_),
    .ZN(_331_));
 NAND2_X1 _798_ (.A1(_326_),
    .A2(_331_),
    .ZN(_332_));
 NAND2_X1 _799_ (.A1(_332_),
    .A2(_174_),
    .ZN(_333_));
 NAND3_X1 _800_ (.A1(_326_),
    .A2(_331_),
    .A3(_135_),
    .ZN(_334_));
 NAND2_X2 _801_ (.A1(_333_),
    .A2(_334_),
    .ZN(resp_msg[15]));
 NAND2_X1 _802_ (.A1(resp_msg[15]),
    .A2(_206_),
    .ZN(_335_));
 NAND2_X1 _803_ (.A1(_322_),
    .A2(_335_),
    .ZN(_336_));
 NAND2_X1 _804_ (.A1(_336_),
    .A2(_186_),
    .ZN(_337_));
 AND2_X1 _805_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .ZN(_338_));
 AOI21_X1 _806_ (.A(_338_),
    .B1(_067_),
    .B2(req_msg[31]),
    .ZN(_339_));
 NAND2_X1 _807_ (.A1(_337_),
    .A2(_339_),
    .ZN(_010_));
 XNOR2_X1 _808_ (.A(_214_),
    .B(_215_),
    .ZN(_340_));
 INV_X1 _809_ (.A(_340_),
    .ZN(resp_msg[1]));
 NAND3_X1 _810_ (.A1(_179_),
    .A2(_181_),
    .A3(resp_msg[1]),
    .ZN(_341_));
 OAI21_X1 _811_ (.A(_341_),
    .B1(_183_),
    .B2(_048_),
    .ZN(_342_));
 NAND2_X1 _812_ (.A1(_342_),
    .A2(_186_),
    .ZN(_343_));
 AND2_X1 _813_ (.A1(_189_),
    .A2(_071_),
    .ZN(_344_));
 AOI21_X1 _814_ (.A(_344_),
    .B1(_067_),
    .B2(req_msg[17]),
    .ZN(_345_));
 NAND2_X1 _815_ (.A1(_343_),
    .A2(_345_),
    .ZN(_011_));
 XNOR2_X1 _816_ (.A(_075_),
    .B(_083_),
    .ZN(resp_msg[2]));
 NAND3_X1 _817_ (.A1(_179_),
    .A2(_181_),
    .A3(resp_msg[2]),
    .ZN(_346_));
 OAI21_X1 _818_ (.A(_346_),
    .B1(_183_),
    .B2(_047_),
    .ZN(_347_));
 NAND2_X1 _819_ (.A1(_347_),
    .A2(_186_),
    .ZN(_348_));
 AND2_X1 _820_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_349_));
 AOI21_X1 _821_ (.A(_349_),
    .B1(_067_),
    .B2(req_msg[18]),
    .ZN(_350_));
 NAND2_X1 _822_ (.A1(_348_),
    .A2(_350_),
    .ZN(_012_));
 XNOR2_X1 _823_ (.A(_220_),
    .B(_079_),
    .ZN(resp_msg[3]));
 NAND3_X1 _824_ (.A1(_179_),
    .A2(_181_),
    .A3(resp_msg[3]),
    .ZN(_351_));
 OAI21_X1 _825_ (.A(_351_),
    .B1(_183_),
    .B2(_046_),
    .ZN(_352_));
 NAND2_X1 _826_ (.A1(_352_),
    .A2(_186_),
    .ZN(_353_));
 AND2_X1 _827_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_354_));
 AOI21_X1 _828_ (.A(_354_),
    .B1(_062_),
    .B2(req_msg[19]),
    .ZN(_355_));
 NAND2_X1 _829_ (.A1(_353_),
    .A2(_355_),
    .ZN(_013_));
 XNOR2_X1 _830_ (.A(_089_),
    .B(_106_),
    .ZN(resp_msg[4]));
 NAND3_X1 _831_ (.A1(_179_),
    .A2(_181_),
    .A3(resp_msg[4]),
    .ZN(_356_));
 OAI21_X1 _832_ (.A(_356_),
    .B1(_183_),
    .B2(_054_),
    .ZN(_357_));
 NAND2_X1 _833_ (.A1(_357_),
    .A2(_185_),
    .ZN(_358_));
 AND2_X1 _834_ (.A1(_188_),
    .A2(\dpath.a_lt_b$in0[4] ),
    .ZN(_359_));
 AOI21_X1 _835_ (.A(_359_),
    .B1(_062_),
    .B2(req_msg[20]),
    .ZN(_360_));
 NAND2_X1 _836_ (.A1(_358_),
    .A2(_360_),
    .ZN(_014_));
 NAND2_X1 _837_ (.A1(_284_),
    .A2(_102_),
    .ZN(_361_));
 INV_X1 _838_ (.A(_102_),
    .ZN(_362_));
 NAND3_X1 _839_ (.A1(_283_),
    .A2(_362_),
    .A3(_231_),
    .ZN(_363_));
 NAND2_X1 _840_ (.A1(_361_),
    .A2(_363_),
    .ZN(resp_msg[5]));
 NAND3_X1 _841_ (.A1(_179_),
    .A2(resp_msg[5]),
    .A3(_181_),
    .ZN(_364_));
 OAI21_X1 _842_ (.A(_364_),
    .B1(_183_),
    .B2(_053_),
    .ZN(_365_));
 NAND2_X1 _843_ (.A1(_365_),
    .A2(_185_),
    .ZN(_366_));
 AND2_X1 _844_ (.A1(_188_),
    .A2(\dpath.a_lt_b$in0[5] ),
    .ZN(_367_));
 AOI21_X1 _845_ (.A(_367_),
    .B1(_062_),
    .B2(req_msg[21]),
    .ZN(_368_));
 NAND2_X1 _846_ (.A1(_366_),
    .A2(_368_),
    .ZN(_015_));
 XNOR2_X1 _847_ (.A(_199_),
    .B(_097_),
    .ZN(resp_msg[6]));
 NAND3_X1 _848_ (.A1(_179_),
    .A2(resp_msg[6]),
    .A3(_181_),
    .ZN(_369_));
 OAI21_X1 _849_ (.A(_369_),
    .B1(_183_),
    .B2(_052_),
    .ZN(_370_));
 NAND2_X1 _850_ (.A1(_370_),
    .A2(_185_),
    .ZN(_371_));
 AND2_X1 _851_ (.A1(_188_),
    .A2(\dpath.a_lt_b$in0[6] ),
    .ZN(_372_));
 AOI21_X1 _852_ (.A(_372_),
    .B1(_062_),
    .B2(req_msg[22]),
    .ZN(_373_));
 NAND2_X1 _853_ (.A1(_371_),
    .A2(_373_),
    .ZN(_016_));
 NAND2_X1 _854_ (.A1(_234_),
    .A2(_093_),
    .ZN(_374_));
 NAND3_X1 _855_ (.A1(_226_),
    .A2(_233_),
    .A3(_238_),
    .ZN(_375_));
 NAND2_X1 _856_ (.A1(_374_),
    .A2(_375_),
    .ZN(resp_msg[7]));
 NAND3_X1 _857_ (.A1(_179_),
    .A2(resp_msg[7]),
    .A3(_181_),
    .ZN(_376_));
 OAI21_X1 _858_ (.A(_376_),
    .B1(_183_),
    .B2(_051_),
    .ZN(_377_));
 NAND2_X1 _859_ (.A1(_377_),
    .A2(_185_),
    .ZN(_378_));
 AND2_X1 _860_ (.A1(_188_),
    .A2(\dpath.a_lt_b$in0[7] ),
    .ZN(_379_));
 AOI21_X1 _861_ (.A(_379_),
    .B1(_062_),
    .B2(req_msg[23]),
    .ZN(_380_));
 NAND2_X1 _862_ (.A1(_378_),
    .A2(_380_),
    .ZN(_017_));
 NAND2_X1 _863_ (.A1(_118_),
    .A2(_156_),
    .ZN(_381_));
 NAND3_X1 _864_ (.A1(_109_),
    .A2(_117_),
    .A3(_157_),
    .ZN(_382_));
 NAND2_X1 _865_ (.A1(_381_),
    .A2(_382_),
    .ZN(resp_msg[8]));
 NAND3_X1 _866_ (.A1(_179_),
    .A2(resp_msg[8]),
    .A3(_181_),
    .ZN(_383_));
 OAI21_X1 _867_ (.A(_383_),
    .B1(_183_),
    .B2(_039_),
    .ZN(_384_));
 NAND2_X1 _868_ (.A1(_384_),
    .A2(_185_),
    .ZN(_385_));
 AND2_X1 _869_ (.A1(_188_),
    .A2(\dpath.a_lt_b$in0[8] ),
    .ZN(_386_));
 AOI21_X1 _870_ (.A(_386_),
    .B1(_062_),
    .B2(req_msg[24]),
    .ZN(_387_));
 NAND2_X1 _871_ (.A1(_385_),
    .A2(_387_),
    .ZN(_018_));
 NAND3_X1 _872_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[9] ),
    .A3(_064_),
    .ZN(_388_));
 NAND2_X1 _873_ (.A1(_213_),
    .A2(_214_),
    .ZN(_389_));
 NOR2_X1 _874_ (.A1(_222_),
    .A2(_389_),
    .ZN(_390_));
 NAND3_X1 _875_ (.A1(_390_),
    .A2(_281_),
    .A3(_215_),
    .ZN(_391_));
 INV_X1 _876_ (.A(_286_),
    .ZN(_392_));
 NAND2_X1 _877_ (.A1(_221_),
    .A2(_218_),
    .ZN(_393_));
 NAND2_X1 _878_ (.A1(_393_),
    .A2(_231_),
    .ZN(_394_));
 NAND2_X1 _879_ (.A1(_394_),
    .A2(_281_),
    .ZN(_395_));
 NAND3_X1 _880_ (.A1(_391_),
    .A2(_392_),
    .A3(_395_),
    .ZN(_396_));
 XNOR2_X1 _881_ (.A(_396_),
    .B(_151_),
    .ZN(resp_msg[9]));
 NAND2_X1 _882_ (.A1(resp_msg[9]),
    .A2(_206_),
    .ZN(_397_));
 NAND2_X1 _883_ (.A1(_388_),
    .A2(_397_),
    .ZN(_398_));
 NAND2_X1 _884_ (.A1(_398_),
    .A2(_185_),
    .ZN(_399_));
 AND2_X1 _885_ (.A1(_188_),
    .A2(\dpath.a_lt_b$in0[9] ),
    .ZN(_400_));
 AOI21_X1 _886_ (.A(_400_),
    .B1(_062_),
    .B2(req_msg[25]),
    .ZN(_401_));
 NAND2_X1 _887_ (.A1(_399_),
    .A2(_401_),
    .ZN(_019_));
 NAND2_X4 _888_ (.A1(_192_),
    .A2(_064_),
    .ZN(_402_));
 BUF_X8 _889_ (.A(_402_),
    .Z(_403_));
 MUX2_X1 _890_ (.A(\dpath.a_lt_b$in0[0] ),
    .B(req_msg[0]),
    .S(_061_),
    .Z(_404_));
 NAND2_X2 _891_ (.A1(_403_),
    .A2(_404_),
    .ZN(_405_));
 BUF_X8 _892_ (.A(_402_),
    .Z(_406_));
 OAI21_X2 _893_ (.A(_405_),
    .B1(_049_),
    .B2(_406_),
    .ZN(_020_));
 NAND2_X1 _894_ (.A1(_066_),
    .A2(req_msg[10]),
    .ZN(_407_));
 OAI21_X1 _895_ (.A(_407_),
    .B1(_062_),
    .B2(_143_),
    .ZN(_408_));
 NAND2_X2 _896_ (.A1(_403_),
    .A2(_408_),
    .ZN(_409_));
 OAI21_X2 _897_ (.A(_409_),
    .B1(_037_),
    .B2(_406_),
    .ZN(_021_));
 NAND2_X1 _898_ (.A1(_066_),
    .A2(req_msg[11]),
    .ZN(_410_));
 OAI21_X1 _899_ (.A(_410_),
    .B1(_062_),
    .B2(_139_),
    .ZN(_411_));
 NAND2_X2 _900_ (.A1(_403_),
    .A2(_411_),
    .ZN(_412_));
 OAI21_X2 _901_ (.A(_412_),
    .B1(_036_),
    .B2(_406_),
    .ZN(_022_));
 NAND2_X1 _902_ (.A1(_066_),
    .A2(req_msg[12]),
    .ZN(_413_));
 CLKBUF_X1 _903_ (.A(_061_),
    .Z(_414_));
 OAI21_X1 _904_ (.A(_413_),
    .B1(_414_),
    .B2(_125_),
    .ZN(_415_));
 NAND2_X2 _905_ (.A1(_403_),
    .A2(_415_),
    .ZN(_416_));
 OAI21_X2 _906_ (.A(_416_),
    .B1(_044_),
    .B2(_406_),
    .ZN(_023_));
 BUF_X8 _907_ (.A(_402_),
    .Z(_417_));
 NAND2_X1 _908_ (.A1(_066_),
    .A2(req_msg[13]),
    .ZN(_418_));
 OAI21_X1 _909_ (.A(_418_),
    .B1(_414_),
    .B2(_119_),
    .ZN(_419_));
 NAND2_X2 _910_ (.A1(_417_),
    .A2(_419_),
    .ZN(_420_));
 OAI21_X2 _911_ (.A(_420_),
    .B1(_043_),
    .B2(_406_),
    .ZN(_024_));
 NAND2_X1 _912_ (.A1(_066_),
    .A2(req_msg[14]),
    .ZN(_421_));
 OAI21_X1 _913_ (.A(_421_),
    .B1(_414_),
    .B2(_131_),
    .ZN(_422_));
 NAND2_X2 _914_ (.A1(_417_),
    .A2(_422_),
    .ZN(_423_));
 OAI21_X2 _915_ (.A(_423_),
    .B1(_042_),
    .B2(_406_),
    .ZN(_025_));
 MUX2_X1 _916_ (.A(\dpath.a_lt_b$in0[15] ),
    .B(req_msg[15]),
    .S(_061_),
    .Z(_424_));
 NAND2_X2 _917_ (.A1(_417_),
    .A2(_424_),
    .ZN(_425_));
 OAI21_X2 _918_ (.A(_425_),
    .B1(_041_),
    .B2(_406_),
    .ZN(_026_));
 MUX2_X1 _919_ (.A(_071_),
    .B(req_msg[1]),
    .S(_061_),
    .Z(_426_));
 NAND2_X2 _920_ (.A1(_417_),
    .A2(_426_),
    .ZN(_427_));
 OAI21_X2 _921_ (.A(_427_),
    .B1(_048_),
    .B2(_406_),
    .ZN(_027_));
 NAND2_X1 _922_ (.A1(_066_),
    .A2(req_msg[2]),
    .ZN(_428_));
 OAI21_X1 _923_ (.A(_428_),
    .B1(_414_),
    .B2(_081_),
    .ZN(_429_));
 NAND2_X2 _924_ (.A1(_417_),
    .A2(_429_),
    .ZN(_430_));
 OAI21_X2 _925_ (.A(_430_),
    .B1(_047_),
    .B2(_406_),
    .ZN(_028_));
 NAND2_X1 _926_ (.A1(_066_),
    .A2(req_msg[3]),
    .ZN(_431_));
 OAI21_X1 _927_ (.A(_431_),
    .B1(_414_),
    .B2(_077_),
    .ZN(_432_));
 NAND2_X2 _928_ (.A1(_417_),
    .A2(_432_),
    .ZN(_433_));
 OAI21_X2 _929_ (.A(_433_),
    .B1(_046_),
    .B2(_406_),
    .ZN(_029_));
 NAND2_X1 _930_ (.A1(_066_),
    .A2(req_msg[4]),
    .ZN(_434_));
 OAI21_X1 _931_ (.A(_434_),
    .B1(_414_),
    .B2(_104_),
    .ZN(_435_));
 NAND2_X2 _932_ (.A1(_417_),
    .A2(_435_),
    .ZN(_436_));
 OAI21_X2 _933_ (.A(_436_),
    .B1(_054_),
    .B2(_403_),
    .ZN(_030_));
 NAND2_X1 _934_ (.A1(_061_),
    .A2(req_msg[5]),
    .ZN(_437_));
 OAI21_X1 _935_ (.A(_437_),
    .B1(_414_),
    .B2(_100_),
    .ZN(_438_));
 NAND2_X2 _936_ (.A1(_417_),
    .A2(_438_),
    .ZN(_439_));
 OAI21_X2 _937_ (.A(_439_),
    .B1(_053_),
    .B2(_403_),
    .ZN(_031_));
 NAND2_X1 _938_ (.A1(_061_),
    .A2(req_msg[6]),
    .ZN(_440_));
 OAI21_X1 _939_ (.A(_440_),
    .B1(_414_),
    .B2(_095_),
    .ZN(_441_));
 NAND2_X2 _940_ (.A1(_417_),
    .A2(_441_),
    .ZN(_442_));
 OAI21_X2 _941_ (.A(_442_),
    .B1(_052_),
    .B2(_403_),
    .ZN(_032_));
 NAND2_X1 _942_ (.A1(_061_),
    .A2(req_msg[7]),
    .ZN(_443_));
 OAI21_X1 _943_ (.A(_443_),
    .B1(_414_),
    .B2(_090_),
    .ZN(_444_));
 NAND2_X2 _944_ (.A1(_417_),
    .A2(_444_),
    .ZN(_445_));
 OAI21_X2 _945_ (.A(_445_),
    .B1(_051_),
    .B2(_403_),
    .ZN(_033_));
 NAND2_X1 _946_ (.A1(_061_),
    .A2(req_msg[8]),
    .ZN(_446_));
 OAI21_X1 _947_ (.A(_446_),
    .B1(_414_),
    .B2(_154_),
    .ZN(_447_));
 NAND2_X1 _948_ (.A1(_402_),
    .A2(_447_),
    .ZN(_448_));
 OAI21_X2 _949_ (.A(_448_),
    .B1(_039_),
    .B2(_403_),
    .ZN(_034_));
 NAND2_X1 _950_ (.A1(_061_),
    .A2(req_msg[9]),
    .ZN(_449_));
 OAI21_X1 _951_ (.A(_449_),
    .B1(_066_),
    .B2(_149_),
    .ZN(_450_));
 NAND2_X1 _952_ (.A1(_402_),
    .A2(_450_),
    .ZN(_451_));
 OAI21_X2 _953_ (.A(_451_),
    .B1(_038_),
    .B2(_403_),
    .ZN(_035_));
 DFF_X1 \ctrl.state.out[0]$_DFF_P_  (.D(_000_),
    .CK(clknet_2_1_0_clk),
    .Q(req_rdy),
    .QN(_003_));
 DFF_X1 \ctrl.state.out[1]$_DFF_P_  (.D(_001_),
    .CK(clknet_2_1_0_clk),
    .Q(\ctrl.state.out[1] ),
    .QN(_485_));
 DFF_X1 \ctrl.state.out[2]$_DFF_P_  (.D(_002_),
    .CK(clknet_2_1_0_clk),
    .Q(\ctrl.state.out[2] ),
    .QN(_484_));
 DFF_X1 \dpath.a_reg.out[0]$_DFFE_PP_  (.D(_004_),
    .CK(clknet_2_3_0_clk),
    .Q(\dpath.a_lt_b$in0[0] ),
    .QN(_483_));
 DFF_X1 \dpath.a_reg.out[10]$_DFFE_PP_  (.D(_005_),
    .CK(clknet_2_0_0_clk),
    .Q(\dpath.a_lt_b$in0[10] ),
    .QN(_482_));
 DFF_X1 \dpath.a_reg.out[11]$_DFFE_PP_  (.D(_006_),
    .CK(clknet_2_2_0_clk),
    .Q(\dpath.a_lt_b$in0[11] ),
    .QN(_481_));
 DFF_X1 \dpath.a_reg.out[12]$_DFFE_PP_  (.D(_007_),
    .CK(clknet_2_0_0_clk),
    .Q(\dpath.a_lt_b$in0[12] ),
    .QN(_480_));
 DFF_X1 \dpath.a_reg.out[13]$_DFFE_PP_  (.D(_008_),
    .CK(clknet_2_2_0_clk),
    .Q(\dpath.a_lt_b$in0[13] ),
    .QN(_479_));
 DFF_X1 \dpath.a_reg.out[14]$_DFFE_PP_  (.D(_009_),
    .CK(clknet_2_0_0_clk),
    .Q(\dpath.a_lt_b$in0[14] ),
    .QN(_478_));
 DFF_X1 \dpath.a_reg.out[15]$_DFFE_PP_  (.D(_010_),
    .CK(clknet_2_0_0_clk),
    .Q(\dpath.a_lt_b$in0[15] ),
    .QN(_477_));
 DFF_X1 \dpath.a_reg.out[1]$_DFFE_PP_  (.D(_011_),
    .CK(clknet_2_0_0_clk),
    .Q(\dpath.a_lt_b$in0[1] ),
    .QN(_476_));
 DFF_X1 \dpath.a_reg.out[2]$_DFFE_PP_  (.D(_012_),
    .CK(clknet_2_2_0_clk),
    .Q(\dpath.a_lt_b$in0[2] ),
    .QN(_475_));
 DFF_X1 \dpath.a_reg.out[3]$_DFFE_PP_  (.D(_013_),
    .CK(clknet_2_2_0_clk),
    .Q(\dpath.a_lt_b$in0[3] ),
    .QN(_474_));
 DFF_X1 \dpath.a_reg.out[4]$_DFFE_PP_  (.D(_014_),
    .CK(clknet_2_3_0_clk),
    .Q(\dpath.a_lt_b$in0[4] ),
    .QN(_473_));
 DFF_X1 \dpath.a_reg.out[5]$_DFFE_PP_  (.D(_015_),
    .CK(clknet_2_3_0_clk),
    .Q(\dpath.a_lt_b$in0[5] ),
    .QN(_472_));
 DFF_X1 \dpath.a_reg.out[6]$_DFFE_PP_  (.D(_016_),
    .CK(clknet_2_3_0_clk),
    .Q(\dpath.a_lt_b$in0[6] ),
    .QN(_471_));
 DFF_X1 \dpath.a_reg.out[7]$_DFFE_PP_  (.D(_017_),
    .CK(clknet_2_1_0_clk),
    .Q(\dpath.a_lt_b$in0[7] ),
    .QN(_470_));
 DFF_X1 \dpath.a_reg.out[8]$_DFFE_PP_  (.D(_018_),
    .CK(clknet_2_1_0_clk),
    .Q(\dpath.a_lt_b$in0[8] ),
    .QN(_469_));
 DFF_X1 \dpath.a_reg.out[9]$_DFFE_PP_  (.D(_019_),
    .CK(clknet_2_3_0_clk),
    .Q(\dpath.a_lt_b$in0[9] ),
    .QN(_468_));
 DFF_X1 \dpath.b_reg.out[0]$_DFFE_PP_  (.D(_020_),
    .CK(clknet_2_3_0_clk),
    .Q(\dpath.a_lt_b$in1[0] ),
    .QN(_467_));
 DFF_X1 \dpath.b_reg.out[10]$_DFFE_PP_  (.D(_021_),
    .CK(clknet_2_2_0_clk),
    .Q(\dpath.a_lt_b$in1[10] ),
    .QN(_466_));
 DFF_X1 \dpath.b_reg.out[11]$_DFFE_PP_  (.D(_022_),
    .CK(clknet_2_2_0_clk),
    .Q(\dpath.a_lt_b$in1[11] ),
    .QN(_465_));
 DFF_X1 \dpath.b_reg.out[12]$_DFFE_PP_  (.D(_023_),
    .CK(clknet_2_0_0_clk),
    .Q(\dpath.a_lt_b$in1[12] ),
    .QN(_464_));
 DFF_X1 \dpath.b_reg.out[13]$_DFFE_PP_  (.D(_024_),
    .CK(clknet_2_2_0_clk),
    .Q(\dpath.a_lt_b$in1[13] ),
    .QN(_463_));
 DFF_X1 \dpath.b_reg.out[14]$_DFFE_PP_  (.D(_025_),
    .CK(clknet_2_0_0_clk),
    .Q(\dpath.a_lt_b$in1[14] ),
    .QN(_462_));
 DFF_X1 \dpath.b_reg.out[15]$_DFFE_PP_  (.D(_026_),
    .CK(clknet_2_0_0_clk),
    .Q(\dpath.a_lt_b$in1[15] ),
    .QN(_461_));
 DFF_X1 \dpath.b_reg.out[1]$_DFFE_PP_  (.D(_027_),
    .CK(clknet_2_1_0_clk),
    .Q(\dpath.a_lt_b$in1[1] ),
    .QN(_460_));
 DFF_X1 \dpath.b_reg.out[2]$_DFFE_PP_  (.D(_028_),
    .CK(clknet_2_2_0_clk),
    .Q(\dpath.a_lt_b$in1[2] ),
    .QN(_459_));
 DFF_X1 \dpath.b_reg.out[3]$_DFFE_PP_  (.D(_029_),
    .CK(clknet_2_2_0_clk),
    .Q(\dpath.a_lt_b$in1[3] ),
    .QN(_458_));
 DFF_X1 \dpath.b_reg.out[4]$_DFFE_PP_  (.D(_030_),
    .CK(clknet_2_3_0_clk),
    .Q(\dpath.a_lt_b$in1[4] ),
    .QN(_457_));
 DFF_X1 \dpath.b_reg.out[5]$_DFFE_PP_  (.D(_031_),
    .CK(clknet_2_3_0_clk),
    .Q(\dpath.a_lt_b$in1[5] ),
    .QN(_456_));
 DFF_X1 \dpath.b_reg.out[6]$_DFFE_PP_  (.D(_032_),
    .CK(clknet_2_3_0_clk),
    .Q(\dpath.a_lt_b$in1[6] ),
    .QN(_455_));
 DFF_X1 \dpath.b_reg.out[7]$_DFFE_PP_  (.D(_033_),
    .CK(clknet_2_1_0_clk),
    .Q(\dpath.a_lt_b$in1[7] ),
    .QN(_454_));
 DFF_X1 \dpath.b_reg.out[8]$_DFFE_PP_  (.D(_034_),
    .CK(clknet_2_1_0_clk),
    .Q(\dpath.a_lt_b$in1[8] ),
    .QN(_453_));
 DFF_X1 \dpath.b_reg.out[9]$_DFFE_PP_  (.D(_035_),
    .CK(clknet_2_3_0_clk),
    .Q(\dpath.a_lt_b$in1[9] ),
    .QN(_452_));
 BUF_X2 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X2 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_0_0_clk));
 BUF_X2 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_1_0_clk));
 BUF_X2 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_2_0_clk));
 BUF_X2 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_3_0_clk));
 BUF_X2 clkload0 (.A(clknet_2_0_0_clk));
 BUF_X2 clkload1 (.A(clknet_2_1_0_clk));
 INV_X1 clkload2 (.A(clknet_2_2_0_clk));
 FILLCELL_X32 FILLCELL_0_0 ();
 FILLCELL_X32 FILLCELL_0_32 ();
 FILLCELL_X32 FILLCELL_0_64 ();
 FILLCELL_X32 FILLCELL_0_96 ();
 FILLCELL_X32 FILLCELL_0_128 ();
 FILLCELL_X32 FILLCELL_0_160 ();
 FILLCELL_X32 FILLCELL_0_192 ();
 FILLCELL_X32 FILLCELL_0_224 ();
 FILLCELL_X32 FILLCELL_0_256 ();
 FILLCELL_X32 FILLCELL_0_288 ();
 FILLCELL_X32 FILLCELL_0_320 ();
 FILLCELL_X32 FILLCELL_0_352 ();
 FILLCELL_X32 FILLCELL_0_384 ();
 FILLCELL_X32 FILLCELL_0_416 ();
 FILLCELL_X32 FILLCELL_0_448 ();
 FILLCELL_X32 FILLCELL_0_480 ();
 FILLCELL_X32 FILLCELL_0_512 ();
 FILLCELL_X32 FILLCELL_0_544 ();
 FILLCELL_X32 FILLCELL_0_576 ();
 FILLCELL_X32 FILLCELL_0_608 ();
 FILLCELL_X32 FILLCELL_0_640 ();
 FILLCELL_X32 FILLCELL_0_672 ();
 FILLCELL_X32 FILLCELL_0_704 ();
 FILLCELL_X32 FILLCELL_0_736 ();
 FILLCELL_X32 FILLCELL_0_768 ();
 FILLCELL_X32 FILLCELL_0_800 ();
 FILLCELL_X32 FILLCELL_0_832 ();
 FILLCELL_X32 FILLCELL_0_864 ();
 FILLCELL_X32 FILLCELL_0_896 ();
 FILLCELL_X32 FILLCELL_0_928 ();
 FILLCELL_X32 FILLCELL_0_960 ();
 FILLCELL_X32 FILLCELL_0_992 ();
 FILLCELL_X32 FILLCELL_0_1024 ();
 FILLCELL_X32 FILLCELL_0_1056 ();
 FILLCELL_X32 FILLCELL_0_1088 ();
 FILLCELL_X32 FILLCELL_0_1120 ();
 FILLCELL_X32 FILLCELL_0_1152 ();
 FILLCELL_X32 FILLCELL_0_1184 ();
 FILLCELL_X32 FILLCELL_0_1216 ();
 FILLCELL_X32 FILLCELL_0_1248 ();
 FILLCELL_X32 FILLCELL_0_1280 ();
 FILLCELL_X32 FILLCELL_0_1312 ();
 FILLCELL_X32 FILLCELL_0_1344 ();
 FILLCELL_X32 FILLCELL_0_1376 ();
 FILLCELL_X32 FILLCELL_0_1408 ();
 FILLCELL_X32 FILLCELL_0_1440 ();
 FILLCELL_X32 FILLCELL_0_1472 ();
 FILLCELL_X32 FILLCELL_0_1504 ();
 FILLCELL_X32 FILLCELL_0_1536 ();
 FILLCELL_X32 FILLCELL_0_1568 ();
 FILLCELL_X32 FILLCELL_0_1600 ();
 FILLCELL_X32 FILLCELL_0_1632 ();
 FILLCELL_X32 FILLCELL_0_1664 ();
 FILLCELL_X32 FILLCELL_0_1696 ();
 FILLCELL_X32 FILLCELL_0_1728 ();
 FILLCELL_X32 FILLCELL_0_1760 ();
 FILLCELL_X32 FILLCELL_0_1792 ();
 FILLCELL_X32 FILLCELL_0_1824 ();
 FILLCELL_X32 FILLCELL_0_1856 ();
 FILLCELL_X8 FILLCELL_0_1888 ();
 FILLCELL_X1 FILLCELL_0_1896 ();
 FILLCELL_X32 FILLCELL_1_0 ();
 FILLCELL_X32 FILLCELL_1_32 ();
 FILLCELL_X32 FILLCELL_1_64 ();
 FILLCELL_X32 FILLCELL_1_96 ();
 FILLCELL_X32 FILLCELL_1_128 ();
 FILLCELL_X32 FILLCELL_1_160 ();
 FILLCELL_X32 FILLCELL_1_192 ();
 FILLCELL_X32 FILLCELL_1_224 ();
 FILLCELL_X32 FILLCELL_1_256 ();
 FILLCELL_X32 FILLCELL_1_288 ();
 FILLCELL_X32 FILLCELL_1_320 ();
 FILLCELL_X32 FILLCELL_1_352 ();
 FILLCELL_X32 FILLCELL_1_384 ();
 FILLCELL_X32 FILLCELL_1_416 ();
 FILLCELL_X32 FILLCELL_1_448 ();
 FILLCELL_X32 FILLCELL_1_480 ();
 FILLCELL_X32 FILLCELL_1_512 ();
 FILLCELL_X32 FILLCELL_1_544 ();
 FILLCELL_X32 FILLCELL_1_576 ();
 FILLCELL_X32 FILLCELL_1_608 ();
 FILLCELL_X32 FILLCELL_1_640 ();
 FILLCELL_X32 FILLCELL_1_672 ();
 FILLCELL_X32 FILLCELL_1_704 ();
 FILLCELL_X32 FILLCELL_1_736 ();
 FILLCELL_X32 FILLCELL_1_768 ();
 FILLCELL_X32 FILLCELL_1_800 ();
 FILLCELL_X32 FILLCELL_1_832 ();
 FILLCELL_X32 FILLCELL_1_864 ();
 FILLCELL_X32 FILLCELL_1_896 ();
 FILLCELL_X32 FILLCELL_1_928 ();
 FILLCELL_X32 FILLCELL_1_960 ();
 FILLCELL_X32 FILLCELL_1_992 ();
 FILLCELL_X32 FILLCELL_1_1024 ();
 FILLCELL_X32 FILLCELL_1_1056 ();
 FILLCELL_X32 FILLCELL_1_1088 ();
 FILLCELL_X32 FILLCELL_1_1120 ();
 FILLCELL_X32 FILLCELL_1_1152 ();
 FILLCELL_X32 FILLCELL_1_1184 ();
 FILLCELL_X32 FILLCELL_1_1216 ();
 FILLCELL_X32 FILLCELL_1_1248 ();
 FILLCELL_X32 FILLCELL_1_1280 ();
 FILLCELL_X32 FILLCELL_1_1312 ();
 FILLCELL_X32 FILLCELL_1_1344 ();
 FILLCELL_X32 FILLCELL_1_1376 ();
 FILLCELL_X32 FILLCELL_1_1408 ();
 FILLCELL_X32 FILLCELL_1_1440 ();
 FILLCELL_X32 FILLCELL_1_1472 ();
 FILLCELL_X32 FILLCELL_1_1504 ();
 FILLCELL_X32 FILLCELL_1_1536 ();
 FILLCELL_X32 FILLCELL_1_1568 ();
 FILLCELL_X32 FILLCELL_1_1600 ();
 FILLCELL_X32 FILLCELL_1_1632 ();
 FILLCELL_X32 FILLCELL_1_1664 ();
 FILLCELL_X32 FILLCELL_1_1696 ();
 FILLCELL_X32 FILLCELL_1_1728 ();
 FILLCELL_X32 FILLCELL_1_1760 ();
 FILLCELL_X32 FILLCELL_1_1792 ();
 FILLCELL_X32 FILLCELL_1_1824 ();
 FILLCELL_X32 FILLCELL_1_1856 ();
 FILLCELL_X8 FILLCELL_1_1888 ();
 FILLCELL_X1 FILLCELL_1_1896 ();
 FILLCELL_X32 FILLCELL_2_0 ();
 FILLCELL_X32 FILLCELL_2_32 ();
 FILLCELL_X32 FILLCELL_2_64 ();
 FILLCELL_X32 FILLCELL_2_96 ();
 FILLCELL_X32 FILLCELL_2_128 ();
 FILLCELL_X32 FILLCELL_2_160 ();
 FILLCELL_X32 FILLCELL_2_192 ();
 FILLCELL_X32 FILLCELL_2_224 ();
 FILLCELL_X32 FILLCELL_2_256 ();
 FILLCELL_X32 FILLCELL_2_288 ();
 FILLCELL_X32 FILLCELL_2_320 ();
 FILLCELL_X32 FILLCELL_2_352 ();
 FILLCELL_X32 FILLCELL_2_384 ();
 FILLCELL_X32 FILLCELL_2_416 ();
 FILLCELL_X32 FILLCELL_2_448 ();
 FILLCELL_X32 FILLCELL_2_480 ();
 FILLCELL_X32 FILLCELL_2_512 ();
 FILLCELL_X32 FILLCELL_2_544 ();
 FILLCELL_X32 FILLCELL_2_576 ();
 FILLCELL_X32 FILLCELL_2_608 ();
 FILLCELL_X32 FILLCELL_2_640 ();
 FILLCELL_X32 FILLCELL_2_672 ();
 FILLCELL_X32 FILLCELL_2_704 ();
 FILLCELL_X32 FILLCELL_2_736 ();
 FILLCELL_X32 FILLCELL_2_768 ();
 FILLCELL_X32 FILLCELL_2_800 ();
 FILLCELL_X32 FILLCELL_2_832 ();
 FILLCELL_X32 FILLCELL_2_864 ();
 FILLCELL_X32 FILLCELL_2_896 ();
 FILLCELL_X32 FILLCELL_2_928 ();
 FILLCELL_X32 FILLCELL_2_960 ();
 FILLCELL_X32 FILLCELL_2_992 ();
 FILLCELL_X32 FILLCELL_2_1024 ();
 FILLCELL_X32 FILLCELL_2_1056 ();
 FILLCELL_X32 FILLCELL_2_1088 ();
 FILLCELL_X32 FILLCELL_2_1120 ();
 FILLCELL_X32 FILLCELL_2_1152 ();
 FILLCELL_X32 FILLCELL_2_1184 ();
 FILLCELL_X32 FILLCELL_2_1216 ();
 FILLCELL_X32 FILLCELL_2_1248 ();
 FILLCELL_X32 FILLCELL_2_1280 ();
 FILLCELL_X32 FILLCELL_2_1312 ();
 FILLCELL_X32 FILLCELL_2_1344 ();
 FILLCELL_X32 FILLCELL_2_1376 ();
 FILLCELL_X32 FILLCELL_2_1408 ();
 FILLCELL_X32 FILLCELL_2_1440 ();
 FILLCELL_X32 FILLCELL_2_1472 ();
 FILLCELL_X32 FILLCELL_2_1504 ();
 FILLCELL_X32 FILLCELL_2_1536 ();
 FILLCELL_X32 FILLCELL_2_1568 ();
 FILLCELL_X32 FILLCELL_2_1600 ();
 FILLCELL_X32 FILLCELL_2_1632 ();
 FILLCELL_X32 FILLCELL_2_1664 ();
 FILLCELL_X32 FILLCELL_2_1696 ();
 FILLCELL_X32 FILLCELL_2_1728 ();
 FILLCELL_X32 FILLCELL_2_1760 ();
 FILLCELL_X32 FILLCELL_2_1792 ();
 FILLCELL_X32 FILLCELL_2_1824 ();
 FILLCELL_X32 FILLCELL_2_1856 ();
 FILLCELL_X8 FILLCELL_2_1888 ();
 FILLCELL_X1 FILLCELL_2_1896 ();
 FILLCELL_X32 FILLCELL_3_0 ();
 FILLCELL_X32 FILLCELL_3_32 ();
 FILLCELL_X32 FILLCELL_3_64 ();
 FILLCELL_X32 FILLCELL_3_96 ();
 FILLCELL_X32 FILLCELL_3_128 ();
 FILLCELL_X32 FILLCELL_3_160 ();
 FILLCELL_X32 FILLCELL_3_192 ();
 FILLCELL_X32 FILLCELL_3_224 ();
 FILLCELL_X32 FILLCELL_3_256 ();
 FILLCELL_X32 FILLCELL_3_288 ();
 FILLCELL_X32 FILLCELL_3_320 ();
 FILLCELL_X32 FILLCELL_3_352 ();
 FILLCELL_X32 FILLCELL_3_384 ();
 FILLCELL_X32 FILLCELL_3_416 ();
 FILLCELL_X32 FILLCELL_3_448 ();
 FILLCELL_X32 FILLCELL_3_480 ();
 FILLCELL_X32 FILLCELL_3_512 ();
 FILLCELL_X32 FILLCELL_3_544 ();
 FILLCELL_X32 FILLCELL_3_576 ();
 FILLCELL_X32 FILLCELL_3_608 ();
 FILLCELL_X32 FILLCELL_3_640 ();
 FILLCELL_X32 FILLCELL_3_672 ();
 FILLCELL_X32 FILLCELL_3_704 ();
 FILLCELL_X32 FILLCELL_3_736 ();
 FILLCELL_X32 FILLCELL_3_768 ();
 FILLCELL_X32 FILLCELL_3_800 ();
 FILLCELL_X32 FILLCELL_3_832 ();
 FILLCELL_X32 FILLCELL_3_864 ();
 FILLCELL_X32 FILLCELL_3_896 ();
 FILLCELL_X32 FILLCELL_3_928 ();
 FILLCELL_X32 FILLCELL_3_960 ();
 FILLCELL_X32 FILLCELL_3_992 ();
 FILLCELL_X32 FILLCELL_3_1024 ();
 FILLCELL_X32 FILLCELL_3_1056 ();
 FILLCELL_X32 FILLCELL_3_1088 ();
 FILLCELL_X32 FILLCELL_3_1120 ();
 FILLCELL_X32 FILLCELL_3_1152 ();
 FILLCELL_X32 FILLCELL_3_1184 ();
 FILLCELL_X32 FILLCELL_3_1216 ();
 FILLCELL_X32 FILLCELL_3_1248 ();
 FILLCELL_X32 FILLCELL_3_1280 ();
 FILLCELL_X32 FILLCELL_3_1312 ();
 FILLCELL_X32 FILLCELL_3_1344 ();
 FILLCELL_X32 FILLCELL_3_1376 ();
 FILLCELL_X32 FILLCELL_3_1408 ();
 FILLCELL_X32 FILLCELL_3_1440 ();
 FILLCELL_X32 FILLCELL_3_1472 ();
 FILLCELL_X32 FILLCELL_3_1504 ();
 FILLCELL_X32 FILLCELL_3_1536 ();
 FILLCELL_X32 FILLCELL_3_1568 ();
 FILLCELL_X32 FILLCELL_3_1600 ();
 FILLCELL_X32 FILLCELL_3_1632 ();
 FILLCELL_X32 FILLCELL_3_1664 ();
 FILLCELL_X32 FILLCELL_3_1696 ();
 FILLCELL_X32 FILLCELL_3_1728 ();
 FILLCELL_X32 FILLCELL_3_1760 ();
 FILLCELL_X32 FILLCELL_3_1792 ();
 FILLCELL_X32 FILLCELL_3_1824 ();
 FILLCELL_X32 FILLCELL_3_1856 ();
 FILLCELL_X8 FILLCELL_3_1888 ();
 FILLCELL_X1 FILLCELL_3_1896 ();
 FILLCELL_X32 FILLCELL_4_0 ();
 FILLCELL_X32 FILLCELL_4_32 ();
 FILLCELL_X32 FILLCELL_4_64 ();
 FILLCELL_X32 FILLCELL_4_96 ();
 FILLCELL_X32 FILLCELL_4_128 ();
 FILLCELL_X32 FILLCELL_4_160 ();
 FILLCELL_X32 FILLCELL_4_192 ();
 FILLCELL_X32 FILLCELL_4_224 ();
 FILLCELL_X32 FILLCELL_4_256 ();
 FILLCELL_X32 FILLCELL_4_288 ();
 FILLCELL_X32 FILLCELL_4_320 ();
 FILLCELL_X32 FILLCELL_4_352 ();
 FILLCELL_X32 FILLCELL_4_384 ();
 FILLCELL_X32 FILLCELL_4_416 ();
 FILLCELL_X32 FILLCELL_4_448 ();
 FILLCELL_X32 FILLCELL_4_480 ();
 FILLCELL_X32 FILLCELL_4_512 ();
 FILLCELL_X32 FILLCELL_4_544 ();
 FILLCELL_X32 FILLCELL_4_576 ();
 FILLCELL_X32 FILLCELL_4_608 ();
 FILLCELL_X32 FILLCELL_4_640 ();
 FILLCELL_X32 FILLCELL_4_672 ();
 FILLCELL_X32 FILLCELL_4_704 ();
 FILLCELL_X32 FILLCELL_4_736 ();
 FILLCELL_X32 FILLCELL_4_768 ();
 FILLCELL_X32 FILLCELL_4_800 ();
 FILLCELL_X32 FILLCELL_4_832 ();
 FILLCELL_X32 FILLCELL_4_864 ();
 FILLCELL_X32 FILLCELL_4_896 ();
 FILLCELL_X32 FILLCELL_4_928 ();
 FILLCELL_X32 FILLCELL_4_960 ();
 FILLCELL_X32 FILLCELL_4_992 ();
 FILLCELL_X32 FILLCELL_4_1024 ();
 FILLCELL_X32 FILLCELL_4_1056 ();
 FILLCELL_X32 FILLCELL_4_1088 ();
 FILLCELL_X32 FILLCELL_4_1120 ();
 FILLCELL_X32 FILLCELL_4_1152 ();
 FILLCELL_X32 FILLCELL_4_1184 ();
 FILLCELL_X32 FILLCELL_4_1216 ();
 FILLCELL_X32 FILLCELL_4_1248 ();
 FILLCELL_X32 FILLCELL_4_1280 ();
 FILLCELL_X32 FILLCELL_4_1312 ();
 FILLCELL_X32 FILLCELL_4_1344 ();
 FILLCELL_X32 FILLCELL_4_1376 ();
 FILLCELL_X32 FILLCELL_4_1408 ();
 FILLCELL_X32 FILLCELL_4_1440 ();
 FILLCELL_X32 FILLCELL_4_1472 ();
 FILLCELL_X32 FILLCELL_4_1504 ();
 FILLCELL_X32 FILLCELL_4_1536 ();
 FILLCELL_X32 FILLCELL_4_1568 ();
 FILLCELL_X32 FILLCELL_4_1600 ();
 FILLCELL_X32 FILLCELL_4_1632 ();
 FILLCELL_X32 FILLCELL_4_1664 ();
 FILLCELL_X32 FILLCELL_4_1696 ();
 FILLCELL_X32 FILLCELL_4_1728 ();
 FILLCELL_X32 FILLCELL_4_1760 ();
 FILLCELL_X32 FILLCELL_4_1792 ();
 FILLCELL_X32 FILLCELL_4_1824 ();
 FILLCELL_X32 FILLCELL_4_1856 ();
 FILLCELL_X8 FILLCELL_4_1888 ();
 FILLCELL_X1 FILLCELL_4_1896 ();
 FILLCELL_X32 FILLCELL_5_0 ();
 FILLCELL_X32 FILLCELL_5_32 ();
 FILLCELL_X32 FILLCELL_5_64 ();
 FILLCELL_X32 FILLCELL_5_96 ();
 FILLCELL_X32 FILLCELL_5_128 ();
 FILLCELL_X32 FILLCELL_5_160 ();
 FILLCELL_X32 FILLCELL_5_192 ();
 FILLCELL_X32 FILLCELL_5_224 ();
 FILLCELL_X32 FILLCELL_5_256 ();
 FILLCELL_X32 FILLCELL_5_288 ();
 FILLCELL_X32 FILLCELL_5_320 ();
 FILLCELL_X32 FILLCELL_5_352 ();
 FILLCELL_X32 FILLCELL_5_384 ();
 FILLCELL_X32 FILLCELL_5_416 ();
 FILLCELL_X32 FILLCELL_5_448 ();
 FILLCELL_X32 FILLCELL_5_480 ();
 FILLCELL_X32 FILLCELL_5_512 ();
 FILLCELL_X32 FILLCELL_5_544 ();
 FILLCELL_X32 FILLCELL_5_576 ();
 FILLCELL_X32 FILLCELL_5_608 ();
 FILLCELL_X32 FILLCELL_5_640 ();
 FILLCELL_X32 FILLCELL_5_672 ();
 FILLCELL_X32 FILLCELL_5_704 ();
 FILLCELL_X32 FILLCELL_5_736 ();
 FILLCELL_X32 FILLCELL_5_768 ();
 FILLCELL_X32 FILLCELL_5_800 ();
 FILLCELL_X32 FILLCELL_5_832 ();
 FILLCELL_X32 FILLCELL_5_864 ();
 FILLCELL_X32 FILLCELL_5_896 ();
 FILLCELL_X32 FILLCELL_5_928 ();
 FILLCELL_X32 FILLCELL_5_960 ();
 FILLCELL_X32 FILLCELL_5_992 ();
 FILLCELL_X32 FILLCELL_5_1024 ();
 FILLCELL_X32 FILLCELL_5_1056 ();
 FILLCELL_X32 FILLCELL_5_1088 ();
 FILLCELL_X32 FILLCELL_5_1120 ();
 FILLCELL_X32 FILLCELL_5_1152 ();
 FILLCELL_X32 FILLCELL_5_1184 ();
 FILLCELL_X32 FILLCELL_5_1216 ();
 FILLCELL_X32 FILLCELL_5_1248 ();
 FILLCELL_X32 FILLCELL_5_1280 ();
 FILLCELL_X32 FILLCELL_5_1312 ();
 FILLCELL_X32 FILLCELL_5_1344 ();
 FILLCELL_X32 FILLCELL_5_1376 ();
 FILLCELL_X32 FILLCELL_5_1408 ();
 FILLCELL_X32 FILLCELL_5_1440 ();
 FILLCELL_X32 FILLCELL_5_1472 ();
 FILLCELL_X32 FILLCELL_5_1504 ();
 FILLCELL_X32 FILLCELL_5_1536 ();
 FILLCELL_X32 FILLCELL_5_1568 ();
 FILLCELL_X32 FILLCELL_5_1600 ();
 FILLCELL_X32 FILLCELL_5_1632 ();
 FILLCELL_X32 FILLCELL_5_1664 ();
 FILLCELL_X32 FILLCELL_5_1696 ();
 FILLCELL_X32 FILLCELL_5_1728 ();
 FILLCELL_X32 FILLCELL_5_1760 ();
 FILLCELL_X32 FILLCELL_5_1792 ();
 FILLCELL_X32 FILLCELL_5_1824 ();
 FILLCELL_X32 FILLCELL_5_1856 ();
 FILLCELL_X8 FILLCELL_5_1888 ();
 FILLCELL_X1 FILLCELL_5_1896 ();
 FILLCELL_X32 FILLCELL_6_0 ();
 FILLCELL_X32 FILLCELL_6_32 ();
 FILLCELL_X32 FILLCELL_6_64 ();
 FILLCELL_X32 FILLCELL_6_96 ();
 FILLCELL_X32 FILLCELL_6_128 ();
 FILLCELL_X32 FILLCELL_6_160 ();
 FILLCELL_X32 FILLCELL_6_192 ();
 FILLCELL_X32 FILLCELL_6_224 ();
 FILLCELL_X32 FILLCELL_6_256 ();
 FILLCELL_X32 FILLCELL_6_288 ();
 FILLCELL_X32 FILLCELL_6_320 ();
 FILLCELL_X32 FILLCELL_6_352 ();
 FILLCELL_X32 FILLCELL_6_384 ();
 FILLCELL_X32 FILLCELL_6_416 ();
 FILLCELL_X32 FILLCELL_6_448 ();
 FILLCELL_X32 FILLCELL_6_480 ();
 FILLCELL_X32 FILLCELL_6_512 ();
 FILLCELL_X32 FILLCELL_6_544 ();
 FILLCELL_X32 FILLCELL_6_576 ();
 FILLCELL_X32 FILLCELL_6_608 ();
 FILLCELL_X32 FILLCELL_6_640 ();
 FILLCELL_X32 FILLCELL_6_672 ();
 FILLCELL_X32 FILLCELL_6_704 ();
 FILLCELL_X32 FILLCELL_6_736 ();
 FILLCELL_X32 FILLCELL_6_768 ();
 FILLCELL_X32 FILLCELL_6_800 ();
 FILLCELL_X32 FILLCELL_6_832 ();
 FILLCELL_X32 FILLCELL_6_864 ();
 FILLCELL_X32 FILLCELL_6_896 ();
 FILLCELL_X32 FILLCELL_6_928 ();
 FILLCELL_X32 FILLCELL_6_960 ();
 FILLCELL_X32 FILLCELL_6_992 ();
 FILLCELL_X32 FILLCELL_6_1024 ();
 FILLCELL_X32 FILLCELL_6_1056 ();
 FILLCELL_X32 FILLCELL_6_1088 ();
 FILLCELL_X32 FILLCELL_6_1120 ();
 FILLCELL_X32 FILLCELL_6_1152 ();
 FILLCELL_X32 FILLCELL_6_1184 ();
 FILLCELL_X32 FILLCELL_6_1216 ();
 FILLCELL_X32 FILLCELL_6_1248 ();
 FILLCELL_X32 FILLCELL_6_1280 ();
 FILLCELL_X32 FILLCELL_6_1312 ();
 FILLCELL_X32 FILLCELL_6_1344 ();
 FILLCELL_X32 FILLCELL_6_1376 ();
 FILLCELL_X32 FILLCELL_6_1408 ();
 FILLCELL_X32 FILLCELL_6_1440 ();
 FILLCELL_X32 FILLCELL_6_1472 ();
 FILLCELL_X32 FILLCELL_6_1504 ();
 FILLCELL_X32 FILLCELL_6_1536 ();
 FILLCELL_X32 FILLCELL_6_1568 ();
 FILLCELL_X32 FILLCELL_6_1600 ();
 FILLCELL_X32 FILLCELL_6_1632 ();
 FILLCELL_X32 FILLCELL_6_1664 ();
 FILLCELL_X32 FILLCELL_6_1696 ();
 FILLCELL_X32 FILLCELL_6_1728 ();
 FILLCELL_X32 FILLCELL_6_1760 ();
 FILLCELL_X32 FILLCELL_6_1792 ();
 FILLCELL_X32 FILLCELL_6_1824 ();
 FILLCELL_X32 FILLCELL_6_1856 ();
 FILLCELL_X8 FILLCELL_6_1888 ();
 FILLCELL_X1 FILLCELL_6_1896 ();
 FILLCELL_X32 FILLCELL_7_0 ();
 FILLCELL_X32 FILLCELL_7_32 ();
 FILLCELL_X32 FILLCELL_7_64 ();
 FILLCELL_X32 FILLCELL_7_96 ();
 FILLCELL_X32 FILLCELL_7_128 ();
 FILLCELL_X32 FILLCELL_7_160 ();
 FILLCELL_X32 FILLCELL_7_192 ();
 FILLCELL_X32 FILLCELL_7_224 ();
 FILLCELL_X32 FILLCELL_7_256 ();
 FILLCELL_X32 FILLCELL_7_288 ();
 FILLCELL_X32 FILLCELL_7_320 ();
 FILLCELL_X32 FILLCELL_7_352 ();
 FILLCELL_X32 FILLCELL_7_384 ();
 FILLCELL_X32 FILLCELL_7_416 ();
 FILLCELL_X32 FILLCELL_7_448 ();
 FILLCELL_X32 FILLCELL_7_480 ();
 FILLCELL_X32 FILLCELL_7_512 ();
 FILLCELL_X32 FILLCELL_7_544 ();
 FILLCELL_X32 FILLCELL_7_576 ();
 FILLCELL_X32 FILLCELL_7_608 ();
 FILLCELL_X32 FILLCELL_7_640 ();
 FILLCELL_X32 FILLCELL_7_672 ();
 FILLCELL_X32 FILLCELL_7_704 ();
 FILLCELL_X32 FILLCELL_7_736 ();
 FILLCELL_X32 FILLCELL_7_768 ();
 FILLCELL_X32 FILLCELL_7_800 ();
 FILLCELL_X32 FILLCELL_7_832 ();
 FILLCELL_X32 FILLCELL_7_864 ();
 FILLCELL_X32 FILLCELL_7_896 ();
 FILLCELL_X32 FILLCELL_7_928 ();
 FILLCELL_X32 FILLCELL_7_960 ();
 FILLCELL_X32 FILLCELL_7_992 ();
 FILLCELL_X32 FILLCELL_7_1024 ();
 FILLCELL_X32 FILLCELL_7_1056 ();
 FILLCELL_X32 FILLCELL_7_1088 ();
 FILLCELL_X32 FILLCELL_7_1120 ();
 FILLCELL_X32 FILLCELL_7_1152 ();
 FILLCELL_X32 FILLCELL_7_1184 ();
 FILLCELL_X32 FILLCELL_7_1216 ();
 FILLCELL_X32 FILLCELL_7_1248 ();
 FILLCELL_X32 FILLCELL_7_1280 ();
 FILLCELL_X32 FILLCELL_7_1312 ();
 FILLCELL_X32 FILLCELL_7_1344 ();
 FILLCELL_X32 FILLCELL_7_1376 ();
 FILLCELL_X32 FILLCELL_7_1408 ();
 FILLCELL_X32 FILLCELL_7_1440 ();
 FILLCELL_X32 FILLCELL_7_1472 ();
 FILLCELL_X32 FILLCELL_7_1504 ();
 FILLCELL_X32 FILLCELL_7_1536 ();
 FILLCELL_X32 FILLCELL_7_1568 ();
 FILLCELL_X32 FILLCELL_7_1600 ();
 FILLCELL_X32 FILLCELL_7_1632 ();
 FILLCELL_X32 FILLCELL_7_1664 ();
 FILLCELL_X32 FILLCELL_7_1696 ();
 FILLCELL_X32 FILLCELL_7_1728 ();
 FILLCELL_X32 FILLCELL_7_1760 ();
 FILLCELL_X32 FILLCELL_7_1792 ();
 FILLCELL_X32 FILLCELL_7_1824 ();
 FILLCELL_X32 FILLCELL_7_1856 ();
 FILLCELL_X8 FILLCELL_7_1888 ();
 FILLCELL_X1 FILLCELL_7_1896 ();
 FILLCELL_X32 FILLCELL_8_0 ();
 FILLCELL_X32 FILLCELL_8_32 ();
 FILLCELL_X32 FILLCELL_8_64 ();
 FILLCELL_X32 FILLCELL_8_96 ();
 FILLCELL_X32 FILLCELL_8_128 ();
 FILLCELL_X32 FILLCELL_8_160 ();
 FILLCELL_X32 FILLCELL_8_192 ();
 FILLCELL_X32 FILLCELL_8_224 ();
 FILLCELL_X32 FILLCELL_8_256 ();
 FILLCELL_X32 FILLCELL_8_288 ();
 FILLCELL_X32 FILLCELL_8_320 ();
 FILLCELL_X32 FILLCELL_8_352 ();
 FILLCELL_X32 FILLCELL_8_384 ();
 FILLCELL_X32 FILLCELL_8_416 ();
 FILLCELL_X32 FILLCELL_8_448 ();
 FILLCELL_X32 FILLCELL_8_480 ();
 FILLCELL_X32 FILLCELL_8_512 ();
 FILLCELL_X32 FILLCELL_8_544 ();
 FILLCELL_X32 FILLCELL_8_576 ();
 FILLCELL_X32 FILLCELL_8_608 ();
 FILLCELL_X32 FILLCELL_8_640 ();
 FILLCELL_X32 FILLCELL_8_672 ();
 FILLCELL_X32 FILLCELL_8_704 ();
 FILLCELL_X32 FILLCELL_8_736 ();
 FILLCELL_X32 FILLCELL_8_768 ();
 FILLCELL_X32 FILLCELL_8_800 ();
 FILLCELL_X32 FILLCELL_8_832 ();
 FILLCELL_X32 FILLCELL_8_864 ();
 FILLCELL_X32 FILLCELL_8_896 ();
 FILLCELL_X32 FILLCELL_8_928 ();
 FILLCELL_X32 FILLCELL_8_960 ();
 FILLCELL_X32 FILLCELL_8_992 ();
 FILLCELL_X32 FILLCELL_8_1024 ();
 FILLCELL_X32 FILLCELL_8_1056 ();
 FILLCELL_X32 FILLCELL_8_1088 ();
 FILLCELL_X32 FILLCELL_8_1120 ();
 FILLCELL_X32 FILLCELL_8_1152 ();
 FILLCELL_X32 FILLCELL_8_1184 ();
 FILLCELL_X32 FILLCELL_8_1216 ();
 FILLCELL_X32 FILLCELL_8_1248 ();
 FILLCELL_X32 FILLCELL_8_1280 ();
 FILLCELL_X32 FILLCELL_8_1312 ();
 FILLCELL_X32 FILLCELL_8_1344 ();
 FILLCELL_X32 FILLCELL_8_1376 ();
 FILLCELL_X32 FILLCELL_8_1408 ();
 FILLCELL_X32 FILLCELL_8_1440 ();
 FILLCELL_X32 FILLCELL_8_1472 ();
 FILLCELL_X32 FILLCELL_8_1504 ();
 FILLCELL_X32 FILLCELL_8_1536 ();
 FILLCELL_X32 FILLCELL_8_1568 ();
 FILLCELL_X32 FILLCELL_8_1600 ();
 FILLCELL_X32 FILLCELL_8_1632 ();
 FILLCELL_X32 FILLCELL_8_1664 ();
 FILLCELL_X32 FILLCELL_8_1696 ();
 FILLCELL_X32 FILLCELL_8_1728 ();
 FILLCELL_X32 FILLCELL_8_1760 ();
 FILLCELL_X32 FILLCELL_8_1792 ();
 FILLCELL_X32 FILLCELL_8_1824 ();
 FILLCELL_X32 FILLCELL_8_1856 ();
 FILLCELL_X8 FILLCELL_8_1888 ();
 FILLCELL_X1 FILLCELL_8_1896 ();
 FILLCELL_X32 FILLCELL_9_0 ();
 FILLCELL_X32 FILLCELL_9_32 ();
 FILLCELL_X32 FILLCELL_9_64 ();
 FILLCELL_X32 FILLCELL_9_96 ();
 FILLCELL_X32 FILLCELL_9_128 ();
 FILLCELL_X32 FILLCELL_9_160 ();
 FILLCELL_X32 FILLCELL_9_192 ();
 FILLCELL_X32 FILLCELL_9_224 ();
 FILLCELL_X32 FILLCELL_9_256 ();
 FILLCELL_X32 FILLCELL_9_288 ();
 FILLCELL_X32 FILLCELL_9_320 ();
 FILLCELL_X32 FILLCELL_9_352 ();
 FILLCELL_X32 FILLCELL_9_384 ();
 FILLCELL_X32 FILLCELL_9_416 ();
 FILLCELL_X32 FILLCELL_9_448 ();
 FILLCELL_X32 FILLCELL_9_480 ();
 FILLCELL_X32 FILLCELL_9_512 ();
 FILLCELL_X32 FILLCELL_9_544 ();
 FILLCELL_X32 FILLCELL_9_576 ();
 FILLCELL_X32 FILLCELL_9_608 ();
 FILLCELL_X32 FILLCELL_9_640 ();
 FILLCELL_X32 FILLCELL_9_672 ();
 FILLCELL_X32 FILLCELL_9_704 ();
 FILLCELL_X32 FILLCELL_9_736 ();
 FILLCELL_X32 FILLCELL_9_768 ();
 FILLCELL_X32 FILLCELL_9_800 ();
 FILLCELL_X32 FILLCELL_9_832 ();
 FILLCELL_X32 FILLCELL_9_864 ();
 FILLCELL_X32 FILLCELL_9_896 ();
 FILLCELL_X32 FILLCELL_9_928 ();
 FILLCELL_X32 FILLCELL_9_960 ();
 FILLCELL_X32 FILLCELL_9_992 ();
 FILLCELL_X32 FILLCELL_9_1024 ();
 FILLCELL_X32 FILLCELL_9_1056 ();
 FILLCELL_X32 FILLCELL_9_1088 ();
 FILLCELL_X32 FILLCELL_9_1120 ();
 FILLCELL_X32 FILLCELL_9_1152 ();
 FILLCELL_X32 FILLCELL_9_1184 ();
 FILLCELL_X32 FILLCELL_9_1216 ();
 FILLCELL_X32 FILLCELL_9_1248 ();
 FILLCELL_X32 FILLCELL_9_1280 ();
 FILLCELL_X32 FILLCELL_9_1312 ();
 FILLCELL_X32 FILLCELL_9_1344 ();
 FILLCELL_X32 FILLCELL_9_1376 ();
 FILLCELL_X32 FILLCELL_9_1408 ();
 FILLCELL_X32 FILLCELL_9_1440 ();
 FILLCELL_X32 FILLCELL_9_1472 ();
 FILLCELL_X32 FILLCELL_9_1504 ();
 FILLCELL_X32 FILLCELL_9_1536 ();
 FILLCELL_X32 FILLCELL_9_1568 ();
 FILLCELL_X32 FILLCELL_9_1600 ();
 FILLCELL_X32 FILLCELL_9_1632 ();
 FILLCELL_X32 FILLCELL_9_1664 ();
 FILLCELL_X32 FILLCELL_9_1696 ();
 FILLCELL_X32 FILLCELL_9_1728 ();
 FILLCELL_X32 FILLCELL_9_1760 ();
 FILLCELL_X32 FILLCELL_9_1792 ();
 FILLCELL_X32 FILLCELL_9_1824 ();
 FILLCELL_X32 FILLCELL_9_1856 ();
 FILLCELL_X8 FILLCELL_9_1888 ();
 FILLCELL_X1 FILLCELL_9_1896 ();
 FILLCELL_X32 FILLCELL_10_0 ();
 FILLCELL_X32 FILLCELL_10_32 ();
 FILLCELL_X32 FILLCELL_10_64 ();
 FILLCELL_X32 FILLCELL_10_96 ();
 FILLCELL_X32 FILLCELL_10_128 ();
 FILLCELL_X32 FILLCELL_10_160 ();
 FILLCELL_X32 FILLCELL_10_192 ();
 FILLCELL_X32 FILLCELL_10_224 ();
 FILLCELL_X32 FILLCELL_10_256 ();
 FILLCELL_X32 FILLCELL_10_288 ();
 FILLCELL_X32 FILLCELL_10_320 ();
 FILLCELL_X32 FILLCELL_10_352 ();
 FILLCELL_X32 FILLCELL_10_384 ();
 FILLCELL_X32 FILLCELL_10_416 ();
 FILLCELL_X32 FILLCELL_10_448 ();
 FILLCELL_X32 FILLCELL_10_480 ();
 FILLCELL_X32 FILLCELL_10_512 ();
 FILLCELL_X32 FILLCELL_10_544 ();
 FILLCELL_X32 FILLCELL_10_576 ();
 FILLCELL_X32 FILLCELL_10_608 ();
 FILLCELL_X32 FILLCELL_10_640 ();
 FILLCELL_X32 FILLCELL_10_672 ();
 FILLCELL_X32 FILLCELL_10_704 ();
 FILLCELL_X32 FILLCELL_10_736 ();
 FILLCELL_X32 FILLCELL_10_768 ();
 FILLCELL_X32 FILLCELL_10_800 ();
 FILLCELL_X32 FILLCELL_10_832 ();
 FILLCELL_X32 FILLCELL_10_864 ();
 FILLCELL_X32 FILLCELL_10_896 ();
 FILLCELL_X32 FILLCELL_10_928 ();
 FILLCELL_X32 FILLCELL_10_960 ();
 FILLCELL_X32 FILLCELL_10_992 ();
 FILLCELL_X32 FILLCELL_10_1024 ();
 FILLCELL_X32 FILLCELL_10_1056 ();
 FILLCELL_X32 FILLCELL_10_1088 ();
 FILLCELL_X32 FILLCELL_10_1120 ();
 FILLCELL_X32 FILLCELL_10_1152 ();
 FILLCELL_X32 FILLCELL_10_1184 ();
 FILLCELL_X32 FILLCELL_10_1216 ();
 FILLCELL_X32 FILLCELL_10_1248 ();
 FILLCELL_X32 FILLCELL_10_1280 ();
 FILLCELL_X32 FILLCELL_10_1312 ();
 FILLCELL_X32 FILLCELL_10_1344 ();
 FILLCELL_X32 FILLCELL_10_1376 ();
 FILLCELL_X32 FILLCELL_10_1408 ();
 FILLCELL_X32 FILLCELL_10_1440 ();
 FILLCELL_X32 FILLCELL_10_1472 ();
 FILLCELL_X32 FILLCELL_10_1504 ();
 FILLCELL_X32 FILLCELL_10_1536 ();
 FILLCELL_X32 FILLCELL_10_1568 ();
 FILLCELL_X32 FILLCELL_10_1600 ();
 FILLCELL_X32 FILLCELL_10_1632 ();
 FILLCELL_X32 FILLCELL_10_1664 ();
 FILLCELL_X32 FILLCELL_10_1696 ();
 FILLCELL_X32 FILLCELL_10_1728 ();
 FILLCELL_X32 FILLCELL_10_1760 ();
 FILLCELL_X32 FILLCELL_10_1792 ();
 FILLCELL_X32 FILLCELL_10_1824 ();
 FILLCELL_X32 FILLCELL_10_1856 ();
 FILLCELL_X8 FILLCELL_10_1888 ();
 FILLCELL_X1 FILLCELL_10_1896 ();
 FILLCELL_X32 FILLCELL_11_0 ();
 FILLCELL_X32 FILLCELL_11_32 ();
 FILLCELL_X32 FILLCELL_11_64 ();
 FILLCELL_X32 FILLCELL_11_96 ();
 FILLCELL_X32 FILLCELL_11_128 ();
 FILLCELL_X32 FILLCELL_11_160 ();
 FILLCELL_X32 FILLCELL_11_192 ();
 FILLCELL_X32 FILLCELL_11_224 ();
 FILLCELL_X32 FILLCELL_11_256 ();
 FILLCELL_X32 FILLCELL_11_288 ();
 FILLCELL_X32 FILLCELL_11_320 ();
 FILLCELL_X32 FILLCELL_11_352 ();
 FILLCELL_X32 FILLCELL_11_384 ();
 FILLCELL_X32 FILLCELL_11_416 ();
 FILLCELL_X32 FILLCELL_11_448 ();
 FILLCELL_X32 FILLCELL_11_480 ();
 FILLCELL_X32 FILLCELL_11_512 ();
 FILLCELL_X32 FILLCELL_11_544 ();
 FILLCELL_X32 FILLCELL_11_576 ();
 FILLCELL_X32 FILLCELL_11_608 ();
 FILLCELL_X32 FILLCELL_11_640 ();
 FILLCELL_X32 FILLCELL_11_672 ();
 FILLCELL_X32 FILLCELL_11_704 ();
 FILLCELL_X32 FILLCELL_11_736 ();
 FILLCELL_X32 FILLCELL_11_768 ();
 FILLCELL_X32 FILLCELL_11_800 ();
 FILLCELL_X32 FILLCELL_11_832 ();
 FILLCELL_X32 FILLCELL_11_864 ();
 FILLCELL_X32 FILLCELL_11_896 ();
 FILLCELL_X32 FILLCELL_11_928 ();
 FILLCELL_X32 FILLCELL_11_960 ();
 FILLCELL_X32 FILLCELL_11_992 ();
 FILLCELL_X32 FILLCELL_11_1024 ();
 FILLCELL_X32 FILLCELL_11_1056 ();
 FILLCELL_X32 FILLCELL_11_1088 ();
 FILLCELL_X32 FILLCELL_11_1120 ();
 FILLCELL_X32 FILLCELL_11_1152 ();
 FILLCELL_X32 FILLCELL_11_1184 ();
 FILLCELL_X32 FILLCELL_11_1216 ();
 FILLCELL_X32 FILLCELL_11_1248 ();
 FILLCELL_X32 FILLCELL_11_1280 ();
 FILLCELL_X32 FILLCELL_11_1312 ();
 FILLCELL_X32 FILLCELL_11_1344 ();
 FILLCELL_X32 FILLCELL_11_1376 ();
 FILLCELL_X32 FILLCELL_11_1408 ();
 FILLCELL_X32 FILLCELL_11_1440 ();
 FILLCELL_X32 FILLCELL_11_1472 ();
 FILLCELL_X32 FILLCELL_11_1504 ();
 FILLCELL_X32 FILLCELL_11_1536 ();
 FILLCELL_X32 FILLCELL_11_1568 ();
 FILLCELL_X32 FILLCELL_11_1600 ();
 FILLCELL_X32 FILLCELL_11_1632 ();
 FILLCELL_X32 FILLCELL_11_1664 ();
 FILLCELL_X32 FILLCELL_11_1696 ();
 FILLCELL_X32 FILLCELL_11_1728 ();
 FILLCELL_X32 FILLCELL_11_1760 ();
 FILLCELL_X32 FILLCELL_11_1792 ();
 FILLCELL_X32 FILLCELL_11_1824 ();
 FILLCELL_X32 FILLCELL_11_1856 ();
 FILLCELL_X8 FILLCELL_11_1888 ();
 FILLCELL_X1 FILLCELL_11_1896 ();
 FILLCELL_X32 FILLCELL_12_0 ();
 FILLCELL_X32 FILLCELL_12_32 ();
 FILLCELL_X32 FILLCELL_12_64 ();
 FILLCELL_X32 FILLCELL_12_96 ();
 FILLCELL_X32 FILLCELL_12_128 ();
 FILLCELL_X32 FILLCELL_12_160 ();
 FILLCELL_X32 FILLCELL_12_192 ();
 FILLCELL_X32 FILLCELL_12_224 ();
 FILLCELL_X32 FILLCELL_12_256 ();
 FILLCELL_X32 FILLCELL_12_288 ();
 FILLCELL_X32 FILLCELL_12_320 ();
 FILLCELL_X32 FILLCELL_12_352 ();
 FILLCELL_X32 FILLCELL_12_384 ();
 FILLCELL_X32 FILLCELL_12_416 ();
 FILLCELL_X32 FILLCELL_12_448 ();
 FILLCELL_X32 FILLCELL_12_480 ();
 FILLCELL_X32 FILLCELL_12_512 ();
 FILLCELL_X32 FILLCELL_12_544 ();
 FILLCELL_X32 FILLCELL_12_576 ();
 FILLCELL_X32 FILLCELL_12_608 ();
 FILLCELL_X32 FILLCELL_12_640 ();
 FILLCELL_X32 FILLCELL_12_672 ();
 FILLCELL_X32 FILLCELL_12_704 ();
 FILLCELL_X32 FILLCELL_12_736 ();
 FILLCELL_X32 FILLCELL_12_768 ();
 FILLCELL_X32 FILLCELL_12_800 ();
 FILLCELL_X32 FILLCELL_12_832 ();
 FILLCELL_X32 FILLCELL_12_864 ();
 FILLCELL_X32 FILLCELL_12_896 ();
 FILLCELL_X32 FILLCELL_12_928 ();
 FILLCELL_X32 FILLCELL_12_960 ();
 FILLCELL_X32 FILLCELL_12_992 ();
 FILLCELL_X32 FILLCELL_12_1024 ();
 FILLCELL_X32 FILLCELL_12_1056 ();
 FILLCELL_X32 FILLCELL_12_1088 ();
 FILLCELL_X32 FILLCELL_12_1120 ();
 FILLCELL_X32 FILLCELL_12_1152 ();
 FILLCELL_X32 FILLCELL_12_1184 ();
 FILLCELL_X32 FILLCELL_12_1216 ();
 FILLCELL_X32 FILLCELL_12_1248 ();
 FILLCELL_X32 FILLCELL_12_1280 ();
 FILLCELL_X32 FILLCELL_12_1312 ();
 FILLCELL_X32 FILLCELL_12_1344 ();
 FILLCELL_X32 FILLCELL_12_1376 ();
 FILLCELL_X32 FILLCELL_12_1408 ();
 FILLCELL_X32 FILLCELL_12_1440 ();
 FILLCELL_X32 FILLCELL_12_1472 ();
 FILLCELL_X32 FILLCELL_12_1504 ();
 FILLCELL_X32 FILLCELL_12_1536 ();
 FILLCELL_X32 FILLCELL_12_1568 ();
 FILLCELL_X32 FILLCELL_12_1600 ();
 FILLCELL_X32 FILLCELL_12_1632 ();
 FILLCELL_X32 FILLCELL_12_1664 ();
 FILLCELL_X32 FILLCELL_12_1696 ();
 FILLCELL_X32 FILLCELL_12_1728 ();
 FILLCELL_X32 FILLCELL_12_1760 ();
 FILLCELL_X32 FILLCELL_12_1792 ();
 FILLCELL_X32 FILLCELL_12_1824 ();
 FILLCELL_X32 FILLCELL_12_1856 ();
 FILLCELL_X8 FILLCELL_12_1888 ();
 FILLCELL_X1 FILLCELL_12_1896 ();
 FILLCELL_X32 FILLCELL_13_0 ();
 FILLCELL_X32 FILLCELL_13_32 ();
 FILLCELL_X32 FILLCELL_13_64 ();
 FILLCELL_X32 FILLCELL_13_96 ();
 FILLCELL_X32 FILLCELL_13_128 ();
 FILLCELL_X32 FILLCELL_13_160 ();
 FILLCELL_X32 FILLCELL_13_192 ();
 FILLCELL_X32 FILLCELL_13_224 ();
 FILLCELL_X32 FILLCELL_13_256 ();
 FILLCELL_X32 FILLCELL_13_288 ();
 FILLCELL_X32 FILLCELL_13_320 ();
 FILLCELL_X32 FILLCELL_13_352 ();
 FILLCELL_X32 FILLCELL_13_384 ();
 FILLCELL_X32 FILLCELL_13_416 ();
 FILLCELL_X32 FILLCELL_13_448 ();
 FILLCELL_X32 FILLCELL_13_480 ();
 FILLCELL_X32 FILLCELL_13_512 ();
 FILLCELL_X32 FILLCELL_13_544 ();
 FILLCELL_X32 FILLCELL_13_576 ();
 FILLCELL_X32 FILLCELL_13_608 ();
 FILLCELL_X32 FILLCELL_13_640 ();
 FILLCELL_X32 FILLCELL_13_672 ();
 FILLCELL_X32 FILLCELL_13_704 ();
 FILLCELL_X32 FILLCELL_13_736 ();
 FILLCELL_X32 FILLCELL_13_768 ();
 FILLCELL_X32 FILLCELL_13_800 ();
 FILLCELL_X32 FILLCELL_13_832 ();
 FILLCELL_X32 FILLCELL_13_864 ();
 FILLCELL_X32 FILLCELL_13_896 ();
 FILLCELL_X32 FILLCELL_13_928 ();
 FILLCELL_X32 FILLCELL_13_960 ();
 FILLCELL_X32 FILLCELL_13_992 ();
 FILLCELL_X32 FILLCELL_13_1024 ();
 FILLCELL_X32 FILLCELL_13_1056 ();
 FILLCELL_X32 FILLCELL_13_1088 ();
 FILLCELL_X32 FILLCELL_13_1120 ();
 FILLCELL_X32 FILLCELL_13_1152 ();
 FILLCELL_X32 FILLCELL_13_1184 ();
 FILLCELL_X32 FILLCELL_13_1216 ();
 FILLCELL_X32 FILLCELL_13_1248 ();
 FILLCELL_X32 FILLCELL_13_1280 ();
 FILLCELL_X32 FILLCELL_13_1312 ();
 FILLCELL_X32 FILLCELL_13_1344 ();
 FILLCELL_X32 FILLCELL_13_1376 ();
 FILLCELL_X32 FILLCELL_13_1408 ();
 FILLCELL_X32 FILLCELL_13_1440 ();
 FILLCELL_X32 FILLCELL_13_1472 ();
 FILLCELL_X32 FILLCELL_13_1504 ();
 FILLCELL_X32 FILLCELL_13_1536 ();
 FILLCELL_X32 FILLCELL_13_1568 ();
 FILLCELL_X32 FILLCELL_13_1600 ();
 FILLCELL_X32 FILLCELL_13_1632 ();
 FILLCELL_X32 FILLCELL_13_1664 ();
 FILLCELL_X32 FILLCELL_13_1696 ();
 FILLCELL_X32 FILLCELL_13_1728 ();
 FILLCELL_X32 FILLCELL_13_1760 ();
 FILLCELL_X32 FILLCELL_13_1792 ();
 FILLCELL_X32 FILLCELL_13_1824 ();
 FILLCELL_X32 FILLCELL_13_1856 ();
 FILLCELL_X8 FILLCELL_13_1888 ();
 FILLCELL_X1 FILLCELL_13_1896 ();
 FILLCELL_X32 FILLCELL_14_0 ();
 FILLCELL_X32 FILLCELL_14_32 ();
 FILLCELL_X32 FILLCELL_14_64 ();
 FILLCELL_X32 FILLCELL_14_96 ();
 FILLCELL_X32 FILLCELL_14_128 ();
 FILLCELL_X32 FILLCELL_14_160 ();
 FILLCELL_X32 FILLCELL_14_192 ();
 FILLCELL_X32 FILLCELL_14_224 ();
 FILLCELL_X32 FILLCELL_14_256 ();
 FILLCELL_X32 FILLCELL_14_288 ();
 FILLCELL_X32 FILLCELL_14_320 ();
 FILLCELL_X32 FILLCELL_14_352 ();
 FILLCELL_X32 FILLCELL_14_384 ();
 FILLCELL_X32 FILLCELL_14_416 ();
 FILLCELL_X32 FILLCELL_14_448 ();
 FILLCELL_X32 FILLCELL_14_480 ();
 FILLCELL_X32 FILLCELL_14_512 ();
 FILLCELL_X32 FILLCELL_14_544 ();
 FILLCELL_X32 FILLCELL_14_576 ();
 FILLCELL_X32 FILLCELL_14_608 ();
 FILLCELL_X32 FILLCELL_14_640 ();
 FILLCELL_X32 FILLCELL_14_672 ();
 FILLCELL_X32 FILLCELL_14_704 ();
 FILLCELL_X32 FILLCELL_14_736 ();
 FILLCELL_X32 FILLCELL_14_768 ();
 FILLCELL_X32 FILLCELL_14_800 ();
 FILLCELL_X32 FILLCELL_14_832 ();
 FILLCELL_X32 FILLCELL_14_864 ();
 FILLCELL_X32 FILLCELL_14_896 ();
 FILLCELL_X32 FILLCELL_14_928 ();
 FILLCELL_X32 FILLCELL_14_960 ();
 FILLCELL_X32 FILLCELL_14_992 ();
 FILLCELL_X32 FILLCELL_14_1024 ();
 FILLCELL_X32 FILLCELL_14_1056 ();
 FILLCELL_X32 FILLCELL_14_1088 ();
 FILLCELL_X32 FILLCELL_14_1120 ();
 FILLCELL_X32 FILLCELL_14_1152 ();
 FILLCELL_X32 FILLCELL_14_1184 ();
 FILLCELL_X32 FILLCELL_14_1216 ();
 FILLCELL_X32 FILLCELL_14_1248 ();
 FILLCELL_X32 FILLCELL_14_1280 ();
 FILLCELL_X32 FILLCELL_14_1312 ();
 FILLCELL_X32 FILLCELL_14_1344 ();
 FILLCELL_X32 FILLCELL_14_1376 ();
 FILLCELL_X32 FILLCELL_14_1408 ();
 FILLCELL_X32 FILLCELL_14_1440 ();
 FILLCELL_X32 FILLCELL_14_1472 ();
 FILLCELL_X32 FILLCELL_14_1504 ();
 FILLCELL_X32 FILLCELL_14_1536 ();
 FILLCELL_X32 FILLCELL_14_1568 ();
 FILLCELL_X32 FILLCELL_14_1600 ();
 FILLCELL_X32 FILLCELL_14_1632 ();
 FILLCELL_X32 FILLCELL_14_1664 ();
 FILLCELL_X32 FILLCELL_14_1696 ();
 FILLCELL_X32 FILLCELL_14_1728 ();
 FILLCELL_X32 FILLCELL_14_1760 ();
 FILLCELL_X32 FILLCELL_14_1792 ();
 FILLCELL_X32 FILLCELL_14_1824 ();
 FILLCELL_X32 FILLCELL_14_1856 ();
 FILLCELL_X8 FILLCELL_14_1888 ();
 FILLCELL_X1 FILLCELL_14_1896 ();
 FILLCELL_X32 FILLCELL_15_0 ();
 FILLCELL_X32 FILLCELL_15_32 ();
 FILLCELL_X32 FILLCELL_15_64 ();
 FILLCELL_X32 FILLCELL_15_96 ();
 FILLCELL_X32 FILLCELL_15_128 ();
 FILLCELL_X32 FILLCELL_15_160 ();
 FILLCELL_X32 FILLCELL_15_192 ();
 FILLCELL_X32 FILLCELL_15_224 ();
 FILLCELL_X32 FILLCELL_15_256 ();
 FILLCELL_X32 FILLCELL_15_288 ();
 FILLCELL_X32 FILLCELL_15_320 ();
 FILLCELL_X32 FILLCELL_15_352 ();
 FILLCELL_X32 FILLCELL_15_384 ();
 FILLCELL_X32 FILLCELL_15_416 ();
 FILLCELL_X32 FILLCELL_15_448 ();
 FILLCELL_X32 FILLCELL_15_480 ();
 FILLCELL_X32 FILLCELL_15_512 ();
 FILLCELL_X32 FILLCELL_15_544 ();
 FILLCELL_X32 FILLCELL_15_576 ();
 FILLCELL_X32 FILLCELL_15_608 ();
 FILLCELL_X32 FILLCELL_15_640 ();
 FILLCELL_X32 FILLCELL_15_672 ();
 FILLCELL_X32 FILLCELL_15_704 ();
 FILLCELL_X32 FILLCELL_15_736 ();
 FILLCELL_X32 FILLCELL_15_768 ();
 FILLCELL_X32 FILLCELL_15_800 ();
 FILLCELL_X32 FILLCELL_15_832 ();
 FILLCELL_X32 FILLCELL_15_864 ();
 FILLCELL_X32 FILLCELL_15_896 ();
 FILLCELL_X32 FILLCELL_15_928 ();
 FILLCELL_X32 FILLCELL_15_960 ();
 FILLCELL_X32 FILLCELL_15_992 ();
 FILLCELL_X32 FILLCELL_15_1024 ();
 FILLCELL_X32 FILLCELL_15_1056 ();
 FILLCELL_X32 FILLCELL_15_1088 ();
 FILLCELL_X32 FILLCELL_15_1120 ();
 FILLCELL_X32 FILLCELL_15_1152 ();
 FILLCELL_X32 FILLCELL_15_1184 ();
 FILLCELL_X32 FILLCELL_15_1216 ();
 FILLCELL_X32 FILLCELL_15_1248 ();
 FILLCELL_X32 FILLCELL_15_1280 ();
 FILLCELL_X32 FILLCELL_15_1312 ();
 FILLCELL_X32 FILLCELL_15_1344 ();
 FILLCELL_X32 FILLCELL_15_1376 ();
 FILLCELL_X32 FILLCELL_15_1408 ();
 FILLCELL_X32 FILLCELL_15_1440 ();
 FILLCELL_X32 FILLCELL_15_1472 ();
 FILLCELL_X32 FILLCELL_15_1504 ();
 FILLCELL_X32 FILLCELL_15_1536 ();
 FILLCELL_X32 FILLCELL_15_1568 ();
 FILLCELL_X32 FILLCELL_15_1600 ();
 FILLCELL_X32 FILLCELL_15_1632 ();
 FILLCELL_X32 FILLCELL_15_1664 ();
 FILLCELL_X32 FILLCELL_15_1696 ();
 FILLCELL_X32 FILLCELL_15_1728 ();
 FILLCELL_X32 FILLCELL_15_1760 ();
 FILLCELL_X32 FILLCELL_15_1792 ();
 FILLCELL_X32 FILLCELL_15_1824 ();
 FILLCELL_X32 FILLCELL_15_1856 ();
 FILLCELL_X8 FILLCELL_15_1888 ();
 FILLCELL_X1 FILLCELL_15_1896 ();
 FILLCELL_X32 FILLCELL_16_0 ();
 FILLCELL_X32 FILLCELL_16_32 ();
 FILLCELL_X32 FILLCELL_16_64 ();
 FILLCELL_X32 FILLCELL_16_96 ();
 FILLCELL_X32 FILLCELL_16_128 ();
 FILLCELL_X32 FILLCELL_16_160 ();
 FILLCELL_X32 FILLCELL_16_192 ();
 FILLCELL_X32 FILLCELL_16_224 ();
 FILLCELL_X32 FILLCELL_16_256 ();
 FILLCELL_X32 FILLCELL_16_288 ();
 FILLCELL_X32 FILLCELL_16_320 ();
 FILLCELL_X32 FILLCELL_16_352 ();
 FILLCELL_X32 FILLCELL_16_384 ();
 FILLCELL_X32 FILLCELL_16_416 ();
 FILLCELL_X32 FILLCELL_16_448 ();
 FILLCELL_X32 FILLCELL_16_480 ();
 FILLCELL_X32 FILLCELL_16_512 ();
 FILLCELL_X32 FILLCELL_16_544 ();
 FILLCELL_X32 FILLCELL_16_576 ();
 FILLCELL_X32 FILLCELL_16_608 ();
 FILLCELL_X32 FILLCELL_16_640 ();
 FILLCELL_X32 FILLCELL_16_672 ();
 FILLCELL_X32 FILLCELL_16_704 ();
 FILLCELL_X32 FILLCELL_16_736 ();
 FILLCELL_X32 FILLCELL_16_768 ();
 FILLCELL_X32 FILLCELL_16_800 ();
 FILLCELL_X32 FILLCELL_16_832 ();
 FILLCELL_X32 FILLCELL_16_864 ();
 FILLCELL_X32 FILLCELL_16_896 ();
 FILLCELL_X32 FILLCELL_16_928 ();
 FILLCELL_X32 FILLCELL_16_960 ();
 FILLCELL_X32 FILLCELL_16_992 ();
 FILLCELL_X32 FILLCELL_16_1024 ();
 FILLCELL_X32 FILLCELL_16_1056 ();
 FILLCELL_X32 FILLCELL_16_1088 ();
 FILLCELL_X32 FILLCELL_16_1120 ();
 FILLCELL_X32 FILLCELL_16_1152 ();
 FILLCELL_X32 FILLCELL_16_1184 ();
 FILLCELL_X32 FILLCELL_16_1216 ();
 FILLCELL_X32 FILLCELL_16_1248 ();
 FILLCELL_X32 FILLCELL_16_1280 ();
 FILLCELL_X32 FILLCELL_16_1312 ();
 FILLCELL_X32 FILLCELL_16_1344 ();
 FILLCELL_X32 FILLCELL_16_1376 ();
 FILLCELL_X32 FILLCELL_16_1408 ();
 FILLCELL_X32 FILLCELL_16_1440 ();
 FILLCELL_X32 FILLCELL_16_1472 ();
 FILLCELL_X32 FILLCELL_16_1504 ();
 FILLCELL_X32 FILLCELL_16_1536 ();
 FILLCELL_X32 FILLCELL_16_1568 ();
 FILLCELL_X32 FILLCELL_16_1600 ();
 FILLCELL_X32 FILLCELL_16_1632 ();
 FILLCELL_X32 FILLCELL_16_1664 ();
 FILLCELL_X32 FILLCELL_16_1696 ();
 FILLCELL_X32 FILLCELL_16_1728 ();
 FILLCELL_X32 FILLCELL_16_1760 ();
 FILLCELL_X32 FILLCELL_16_1792 ();
 FILLCELL_X32 FILLCELL_16_1824 ();
 FILLCELL_X32 FILLCELL_16_1856 ();
 FILLCELL_X8 FILLCELL_16_1888 ();
 FILLCELL_X1 FILLCELL_16_1896 ();
 FILLCELL_X32 FILLCELL_17_0 ();
 FILLCELL_X32 FILLCELL_17_32 ();
 FILLCELL_X32 FILLCELL_17_64 ();
 FILLCELL_X32 FILLCELL_17_96 ();
 FILLCELL_X32 FILLCELL_17_128 ();
 FILLCELL_X32 FILLCELL_17_160 ();
 FILLCELL_X32 FILLCELL_17_192 ();
 FILLCELL_X32 FILLCELL_17_224 ();
 FILLCELL_X32 FILLCELL_17_256 ();
 FILLCELL_X32 FILLCELL_17_288 ();
 FILLCELL_X32 FILLCELL_17_320 ();
 FILLCELL_X32 FILLCELL_17_352 ();
 FILLCELL_X32 FILLCELL_17_384 ();
 FILLCELL_X32 FILLCELL_17_416 ();
 FILLCELL_X32 FILLCELL_17_448 ();
 FILLCELL_X32 FILLCELL_17_480 ();
 FILLCELL_X32 FILLCELL_17_512 ();
 FILLCELL_X32 FILLCELL_17_544 ();
 FILLCELL_X32 FILLCELL_17_576 ();
 FILLCELL_X32 FILLCELL_17_608 ();
 FILLCELL_X32 FILLCELL_17_640 ();
 FILLCELL_X32 FILLCELL_17_672 ();
 FILLCELL_X32 FILLCELL_17_704 ();
 FILLCELL_X32 FILLCELL_17_736 ();
 FILLCELL_X32 FILLCELL_17_768 ();
 FILLCELL_X32 FILLCELL_17_800 ();
 FILLCELL_X32 FILLCELL_17_832 ();
 FILLCELL_X32 FILLCELL_17_864 ();
 FILLCELL_X32 FILLCELL_17_896 ();
 FILLCELL_X32 FILLCELL_17_928 ();
 FILLCELL_X32 FILLCELL_17_960 ();
 FILLCELL_X32 FILLCELL_17_992 ();
 FILLCELL_X32 FILLCELL_17_1024 ();
 FILLCELL_X32 FILLCELL_17_1056 ();
 FILLCELL_X32 FILLCELL_17_1088 ();
 FILLCELL_X32 FILLCELL_17_1120 ();
 FILLCELL_X32 FILLCELL_17_1152 ();
 FILLCELL_X32 FILLCELL_17_1184 ();
 FILLCELL_X32 FILLCELL_17_1216 ();
 FILLCELL_X32 FILLCELL_17_1248 ();
 FILLCELL_X32 FILLCELL_17_1280 ();
 FILLCELL_X32 FILLCELL_17_1312 ();
 FILLCELL_X32 FILLCELL_17_1344 ();
 FILLCELL_X32 FILLCELL_17_1376 ();
 FILLCELL_X32 FILLCELL_17_1408 ();
 FILLCELL_X32 FILLCELL_17_1440 ();
 FILLCELL_X32 FILLCELL_17_1472 ();
 FILLCELL_X32 FILLCELL_17_1504 ();
 FILLCELL_X32 FILLCELL_17_1536 ();
 FILLCELL_X32 FILLCELL_17_1568 ();
 FILLCELL_X32 FILLCELL_17_1600 ();
 FILLCELL_X32 FILLCELL_17_1632 ();
 FILLCELL_X32 FILLCELL_17_1664 ();
 FILLCELL_X32 FILLCELL_17_1696 ();
 FILLCELL_X32 FILLCELL_17_1728 ();
 FILLCELL_X32 FILLCELL_17_1760 ();
 FILLCELL_X32 FILLCELL_17_1792 ();
 FILLCELL_X32 FILLCELL_17_1824 ();
 FILLCELL_X32 FILLCELL_17_1856 ();
 FILLCELL_X8 FILLCELL_17_1888 ();
 FILLCELL_X1 FILLCELL_17_1896 ();
 FILLCELL_X32 FILLCELL_18_0 ();
 FILLCELL_X32 FILLCELL_18_32 ();
 FILLCELL_X32 FILLCELL_18_64 ();
 FILLCELL_X32 FILLCELL_18_96 ();
 FILLCELL_X32 FILLCELL_18_128 ();
 FILLCELL_X32 FILLCELL_18_160 ();
 FILLCELL_X32 FILLCELL_18_192 ();
 FILLCELL_X32 FILLCELL_18_224 ();
 FILLCELL_X32 FILLCELL_18_256 ();
 FILLCELL_X32 FILLCELL_18_288 ();
 FILLCELL_X32 FILLCELL_18_320 ();
 FILLCELL_X32 FILLCELL_18_352 ();
 FILLCELL_X32 FILLCELL_18_384 ();
 FILLCELL_X32 FILLCELL_18_416 ();
 FILLCELL_X32 FILLCELL_18_448 ();
 FILLCELL_X32 FILLCELL_18_480 ();
 FILLCELL_X32 FILLCELL_18_512 ();
 FILLCELL_X32 FILLCELL_18_544 ();
 FILLCELL_X32 FILLCELL_18_576 ();
 FILLCELL_X32 FILLCELL_18_608 ();
 FILLCELL_X32 FILLCELL_18_640 ();
 FILLCELL_X32 FILLCELL_18_672 ();
 FILLCELL_X32 FILLCELL_18_704 ();
 FILLCELL_X32 FILLCELL_18_736 ();
 FILLCELL_X32 FILLCELL_18_768 ();
 FILLCELL_X32 FILLCELL_18_800 ();
 FILLCELL_X32 FILLCELL_18_832 ();
 FILLCELL_X32 FILLCELL_18_864 ();
 FILLCELL_X32 FILLCELL_18_896 ();
 FILLCELL_X32 FILLCELL_18_928 ();
 FILLCELL_X32 FILLCELL_18_960 ();
 FILLCELL_X32 FILLCELL_18_992 ();
 FILLCELL_X32 FILLCELL_18_1024 ();
 FILLCELL_X32 FILLCELL_18_1056 ();
 FILLCELL_X32 FILLCELL_18_1088 ();
 FILLCELL_X32 FILLCELL_18_1120 ();
 FILLCELL_X32 FILLCELL_18_1152 ();
 FILLCELL_X32 FILLCELL_18_1184 ();
 FILLCELL_X32 FILLCELL_18_1216 ();
 FILLCELL_X32 FILLCELL_18_1248 ();
 FILLCELL_X32 FILLCELL_18_1280 ();
 FILLCELL_X32 FILLCELL_18_1312 ();
 FILLCELL_X32 FILLCELL_18_1344 ();
 FILLCELL_X32 FILLCELL_18_1376 ();
 FILLCELL_X32 FILLCELL_18_1408 ();
 FILLCELL_X32 FILLCELL_18_1440 ();
 FILLCELL_X32 FILLCELL_18_1472 ();
 FILLCELL_X32 FILLCELL_18_1504 ();
 FILLCELL_X32 FILLCELL_18_1536 ();
 FILLCELL_X32 FILLCELL_18_1568 ();
 FILLCELL_X32 FILLCELL_18_1600 ();
 FILLCELL_X32 FILLCELL_18_1632 ();
 FILLCELL_X32 FILLCELL_18_1664 ();
 FILLCELL_X32 FILLCELL_18_1696 ();
 FILLCELL_X32 FILLCELL_18_1728 ();
 FILLCELL_X32 FILLCELL_18_1760 ();
 FILLCELL_X32 FILLCELL_18_1792 ();
 FILLCELL_X32 FILLCELL_18_1824 ();
 FILLCELL_X32 FILLCELL_18_1856 ();
 FILLCELL_X8 FILLCELL_18_1888 ();
 FILLCELL_X1 FILLCELL_18_1896 ();
 FILLCELL_X32 FILLCELL_19_0 ();
 FILLCELL_X32 FILLCELL_19_32 ();
 FILLCELL_X32 FILLCELL_19_64 ();
 FILLCELL_X32 FILLCELL_19_96 ();
 FILLCELL_X32 FILLCELL_19_128 ();
 FILLCELL_X32 FILLCELL_19_160 ();
 FILLCELL_X32 FILLCELL_19_192 ();
 FILLCELL_X32 FILLCELL_19_224 ();
 FILLCELL_X32 FILLCELL_19_256 ();
 FILLCELL_X32 FILLCELL_19_288 ();
 FILLCELL_X32 FILLCELL_19_320 ();
 FILLCELL_X32 FILLCELL_19_352 ();
 FILLCELL_X32 FILLCELL_19_384 ();
 FILLCELL_X32 FILLCELL_19_416 ();
 FILLCELL_X32 FILLCELL_19_448 ();
 FILLCELL_X32 FILLCELL_19_480 ();
 FILLCELL_X32 FILLCELL_19_512 ();
 FILLCELL_X32 FILLCELL_19_544 ();
 FILLCELL_X32 FILLCELL_19_576 ();
 FILLCELL_X32 FILLCELL_19_608 ();
 FILLCELL_X32 FILLCELL_19_640 ();
 FILLCELL_X32 FILLCELL_19_672 ();
 FILLCELL_X32 FILLCELL_19_704 ();
 FILLCELL_X32 FILLCELL_19_736 ();
 FILLCELL_X32 FILLCELL_19_768 ();
 FILLCELL_X32 FILLCELL_19_800 ();
 FILLCELL_X32 FILLCELL_19_832 ();
 FILLCELL_X32 FILLCELL_19_864 ();
 FILLCELL_X32 FILLCELL_19_896 ();
 FILLCELL_X32 FILLCELL_19_928 ();
 FILLCELL_X32 FILLCELL_19_960 ();
 FILLCELL_X32 FILLCELL_19_992 ();
 FILLCELL_X32 FILLCELL_19_1024 ();
 FILLCELL_X32 FILLCELL_19_1056 ();
 FILLCELL_X32 FILLCELL_19_1088 ();
 FILLCELL_X32 FILLCELL_19_1120 ();
 FILLCELL_X32 FILLCELL_19_1152 ();
 FILLCELL_X32 FILLCELL_19_1184 ();
 FILLCELL_X32 FILLCELL_19_1216 ();
 FILLCELL_X32 FILLCELL_19_1248 ();
 FILLCELL_X32 FILLCELL_19_1280 ();
 FILLCELL_X32 FILLCELL_19_1312 ();
 FILLCELL_X32 FILLCELL_19_1344 ();
 FILLCELL_X32 FILLCELL_19_1376 ();
 FILLCELL_X32 FILLCELL_19_1408 ();
 FILLCELL_X32 FILLCELL_19_1440 ();
 FILLCELL_X32 FILLCELL_19_1472 ();
 FILLCELL_X32 FILLCELL_19_1504 ();
 FILLCELL_X32 FILLCELL_19_1536 ();
 FILLCELL_X32 FILLCELL_19_1568 ();
 FILLCELL_X32 FILLCELL_19_1600 ();
 FILLCELL_X32 FILLCELL_19_1632 ();
 FILLCELL_X32 FILLCELL_19_1664 ();
 FILLCELL_X32 FILLCELL_19_1696 ();
 FILLCELL_X32 FILLCELL_19_1728 ();
 FILLCELL_X32 FILLCELL_19_1760 ();
 FILLCELL_X32 FILLCELL_19_1792 ();
 FILLCELL_X32 FILLCELL_19_1824 ();
 FILLCELL_X32 FILLCELL_19_1856 ();
 FILLCELL_X8 FILLCELL_19_1888 ();
 FILLCELL_X1 FILLCELL_19_1896 ();
 FILLCELL_X32 FILLCELL_20_0 ();
 FILLCELL_X32 FILLCELL_20_32 ();
 FILLCELL_X32 FILLCELL_20_64 ();
 FILLCELL_X32 FILLCELL_20_96 ();
 FILLCELL_X32 FILLCELL_20_128 ();
 FILLCELL_X32 FILLCELL_20_160 ();
 FILLCELL_X32 FILLCELL_20_192 ();
 FILLCELL_X32 FILLCELL_20_224 ();
 FILLCELL_X32 FILLCELL_20_256 ();
 FILLCELL_X32 FILLCELL_20_288 ();
 FILLCELL_X32 FILLCELL_20_320 ();
 FILLCELL_X32 FILLCELL_20_352 ();
 FILLCELL_X32 FILLCELL_20_384 ();
 FILLCELL_X32 FILLCELL_20_416 ();
 FILLCELL_X32 FILLCELL_20_448 ();
 FILLCELL_X32 FILLCELL_20_480 ();
 FILLCELL_X32 FILLCELL_20_512 ();
 FILLCELL_X32 FILLCELL_20_544 ();
 FILLCELL_X32 FILLCELL_20_576 ();
 FILLCELL_X32 FILLCELL_20_608 ();
 FILLCELL_X32 FILLCELL_20_640 ();
 FILLCELL_X32 FILLCELL_20_672 ();
 FILLCELL_X32 FILLCELL_20_704 ();
 FILLCELL_X32 FILLCELL_20_736 ();
 FILLCELL_X32 FILLCELL_20_768 ();
 FILLCELL_X32 FILLCELL_20_800 ();
 FILLCELL_X32 FILLCELL_20_832 ();
 FILLCELL_X32 FILLCELL_20_864 ();
 FILLCELL_X32 FILLCELL_20_896 ();
 FILLCELL_X32 FILLCELL_20_928 ();
 FILLCELL_X32 FILLCELL_20_960 ();
 FILLCELL_X32 FILLCELL_20_992 ();
 FILLCELL_X32 FILLCELL_20_1024 ();
 FILLCELL_X32 FILLCELL_20_1056 ();
 FILLCELL_X32 FILLCELL_20_1088 ();
 FILLCELL_X32 FILLCELL_20_1120 ();
 FILLCELL_X32 FILLCELL_20_1152 ();
 FILLCELL_X32 FILLCELL_20_1184 ();
 FILLCELL_X32 FILLCELL_20_1216 ();
 FILLCELL_X32 FILLCELL_20_1248 ();
 FILLCELL_X32 FILLCELL_20_1280 ();
 FILLCELL_X32 FILLCELL_20_1312 ();
 FILLCELL_X32 FILLCELL_20_1344 ();
 FILLCELL_X32 FILLCELL_20_1376 ();
 FILLCELL_X32 FILLCELL_20_1408 ();
 FILLCELL_X32 FILLCELL_20_1440 ();
 FILLCELL_X32 FILLCELL_20_1472 ();
 FILLCELL_X32 FILLCELL_20_1504 ();
 FILLCELL_X32 FILLCELL_20_1536 ();
 FILLCELL_X32 FILLCELL_20_1568 ();
 FILLCELL_X32 FILLCELL_20_1600 ();
 FILLCELL_X32 FILLCELL_20_1632 ();
 FILLCELL_X32 FILLCELL_20_1664 ();
 FILLCELL_X32 FILLCELL_20_1696 ();
 FILLCELL_X32 FILLCELL_20_1728 ();
 FILLCELL_X32 FILLCELL_20_1760 ();
 FILLCELL_X32 FILLCELL_20_1792 ();
 FILLCELL_X32 FILLCELL_20_1824 ();
 FILLCELL_X32 FILLCELL_20_1856 ();
 FILLCELL_X8 FILLCELL_20_1888 ();
 FILLCELL_X1 FILLCELL_20_1896 ();
 FILLCELL_X32 FILLCELL_21_0 ();
 FILLCELL_X32 FILLCELL_21_32 ();
 FILLCELL_X32 FILLCELL_21_64 ();
 FILLCELL_X32 FILLCELL_21_96 ();
 FILLCELL_X32 FILLCELL_21_128 ();
 FILLCELL_X32 FILLCELL_21_160 ();
 FILLCELL_X32 FILLCELL_21_192 ();
 FILLCELL_X32 FILLCELL_21_224 ();
 FILLCELL_X32 FILLCELL_21_256 ();
 FILLCELL_X32 FILLCELL_21_288 ();
 FILLCELL_X32 FILLCELL_21_320 ();
 FILLCELL_X32 FILLCELL_21_352 ();
 FILLCELL_X32 FILLCELL_21_384 ();
 FILLCELL_X32 FILLCELL_21_416 ();
 FILLCELL_X32 FILLCELL_21_448 ();
 FILLCELL_X32 FILLCELL_21_480 ();
 FILLCELL_X32 FILLCELL_21_512 ();
 FILLCELL_X32 FILLCELL_21_544 ();
 FILLCELL_X32 FILLCELL_21_576 ();
 FILLCELL_X32 FILLCELL_21_608 ();
 FILLCELL_X32 FILLCELL_21_640 ();
 FILLCELL_X32 FILLCELL_21_672 ();
 FILLCELL_X32 FILLCELL_21_704 ();
 FILLCELL_X32 FILLCELL_21_736 ();
 FILLCELL_X32 FILLCELL_21_768 ();
 FILLCELL_X32 FILLCELL_21_800 ();
 FILLCELL_X32 FILLCELL_21_832 ();
 FILLCELL_X32 FILLCELL_21_864 ();
 FILLCELL_X32 FILLCELL_21_896 ();
 FILLCELL_X32 FILLCELL_21_928 ();
 FILLCELL_X32 FILLCELL_21_960 ();
 FILLCELL_X32 FILLCELL_21_992 ();
 FILLCELL_X32 FILLCELL_21_1024 ();
 FILLCELL_X32 FILLCELL_21_1056 ();
 FILLCELL_X32 FILLCELL_21_1088 ();
 FILLCELL_X32 FILLCELL_21_1120 ();
 FILLCELL_X32 FILLCELL_21_1152 ();
 FILLCELL_X32 FILLCELL_21_1184 ();
 FILLCELL_X32 FILLCELL_21_1216 ();
 FILLCELL_X32 FILLCELL_21_1248 ();
 FILLCELL_X32 FILLCELL_21_1280 ();
 FILLCELL_X32 FILLCELL_21_1312 ();
 FILLCELL_X32 FILLCELL_21_1344 ();
 FILLCELL_X32 FILLCELL_21_1376 ();
 FILLCELL_X32 FILLCELL_21_1408 ();
 FILLCELL_X32 FILLCELL_21_1440 ();
 FILLCELL_X32 FILLCELL_21_1472 ();
 FILLCELL_X32 FILLCELL_21_1504 ();
 FILLCELL_X32 FILLCELL_21_1536 ();
 FILLCELL_X32 FILLCELL_21_1568 ();
 FILLCELL_X32 FILLCELL_21_1600 ();
 FILLCELL_X32 FILLCELL_21_1632 ();
 FILLCELL_X32 FILLCELL_21_1664 ();
 FILLCELL_X32 FILLCELL_21_1696 ();
 FILLCELL_X32 FILLCELL_21_1728 ();
 FILLCELL_X32 FILLCELL_21_1760 ();
 FILLCELL_X32 FILLCELL_21_1792 ();
 FILLCELL_X32 FILLCELL_21_1824 ();
 FILLCELL_X32 FILLCELL_21_1856 ();
 FILLCELL_X8 FILLCELL_21_1888 ();
 FILLCELL_X1 FILLCELL_21_1896 ();
 FILLCELL_X32 FILLCELL_22_0 ();
 FILLCELL_X32 FILLCELL_22_32 ();
 FILLCELL_X32 FILLCELL_22_64 ();
 FILLCELL_X32 FILLCELL_22_96 ();
 FILLCELL_X32 FILLCELL_22_128 ();
 FILLCELL_X32 FILLCELL_22_160 ();
 FILLCELL_X32 FILLCELL_22_192 ();
 FILLCELL_X32 FILLCELL_22_224 ();
 FILLCELL_X32 FILLCELL_22_256 ();
 FILLCELL_X32 FILLCELL_22_288 ();
 FILLCELL_X32 FILLCELL_22_320 ();
 FILLCELL_X32 FILLCELL_22_352 ();
 FILLCELL_X32 FILLCELL_22_384 ();
 FILLCELL_X32 FILLCELL_22_416 ();
 FILLCELL_X32 FILLCELL_22_448 ();
 FILLCELL_X32 FILLCELL_22_480 ();
 FILLCELL_X32 FILLCELL_22_512 ();
 FILLCELL_X32 FILLCELL_22_544 ();
 FILLCELL_X32 FILLCELL_22_576 ();
 FILLCELL_X32 FILLCELL_22_608 ();
 FILLCELL_X32 FILLCELL_22_640 ();
 FILLCELL_X32 FILLCELL_22_672 ();
 FILLCELL_X32 FILLCELL_22_704 ();
 FILLCELL_X32 FILLCELL_22_736 ();
 FILLCELL_X32 FILLCELL_22_768 ();
 FILLCELL_X32 FILLCELL_22_800 ();
 FILLCELL_X32 FILLCELL_22_832 ();
 FILLCELL_X32 FILLCELL_22_864 ();
 FILLCELL_X32 FILLCELL_22_896 ();
 FILLCELL_X32 FILLCELL_22_928 ();
 FILLCELL_X32 FILLCELL_22_960 ();
 FILLCELL_X32 FILLCELL_22_992 ();
 FILLCELL_X32 FILLCELL_22_1024 ();
 FILLCELL_X32 FILLCELL_22_1056 ();
 FILLCELL_X32 FILLCELL_22_1088 ();
 FILLCELL_X32 FILLCELL_22_1120 ();
 FILLCELL_X32 FILLCELL_22_1152 ();
 FILLCELL_X32 FILLCELL_22_1184 ();
 FILLCELL_X32 FILLCELL_22_1216 ();
 FILLCELL_X32 FILLCELL_22_1248 ();
 FILLCELL_X32 FILLCELL_22_1280 ();
 FILLCELL_X32 FILLCELL_22_1312 ();
 FILLCELL_X32 FILLCELL_22_1344 ();
 FILLCELL_X32 FILLCELL_22_1376 ();
 FILLCELL_X32 FILLCELL_22_1408 ();
 FILLCELL_X32 FILLCELL_22_1440 ();
 FILLCELL_X32 FILLCELL_22_1472 ();
 FILLCELL_X32 FILLCELL_22_1504 ();
 FILLCELL_X32 FILLCELL_22_1536 ();
 FILLCELL_X32 FILLCELL_22_1568 ();
 FILLCELL_X32 FILLCELL_22_1600 ();
 FILLCELL_X32 FILLCELL_22_1632 ();
 FILLCELL_X32 FILLCELL_22_1664 ();
 FILLCELL_X32 FILLCELL_22_1696 ();
 FILLCELL_X32 FILLCELL_22_1728 ();
 FILLCELL_X32 FILLCELL_22_1760 ();
 FILLCELL_X32 FILLCELL_22_1792 ();
 FILLCELL_X32 FILLCELL_22_1824 ();
 FILLCELL_X32 FILLCELL_22_1856 ();
 FILLCELL_X8 FILLCELL_22_1888 ();
 FILLCELL_X1 FILLCELL_22_1896 ();
 FILLCELL_X32 FILLCELL_23_0 ();
 FILLCELL_X32 FILLCELL_23_32 ();
 FILLCELL_X32 FILLCELL_23_64 ();
 FILLCELL_X32 FILLCELL_23_96 ();
 FILLCELL_X32 FILLCELL_23_128 ();
 FILLCELL_X32 FILLCELL_23_160 ();
 FILLCELL_X32 FILLCELL_23_192 ();
 FILLCELL_X32 FILLCELL_23_224 ();
 FILLCELL_X32 FILLCELL_23_256 ();
 FILLCELL_X32 FILLCELL_23_288 ();
 FILLCELL_X32 FILLCELL_23_320 ();
 FILLCELL_X32 FILLCELL_23_352 ();
 FILLCELL_X32 FILLCELL_23_384 ();
 FILLCELL_X32 FILLCELL_23_416 ();
 FILLCELL_X32 FILLCELL_23_448 ();
 FILLCELL_X32 FILLCELL_23_480 ();
 FILLCELL_X32 FILLCELL_23_512 ();
 FILLCELL_X32 FILLCELL_23_544 ();
 FILLCELL_X32 FILLCELL_23_576 ();
 FILLCELL_X32 FILLCELL_23_608 ();
 FILLCELL_X32 FILLCELL_23_640 ();
 FILLCELL_X32 FILLCELL_23_672 ();
 FILLCELL_X32 FILLCELL_23_704 ();
 FILLCELL_X32 FILLCELL_23_736 ();
 FILLCELL_X32 FILLCELL_23_768 ();
 FILLCELL_X32 FILLCELL_23_800 ();
 FILLCELL_X32 FILLCELL_23_832 ();
 FILLCELL_X32 FILLCELL_23_864 ();
 FILLCELL_X32 FILLCELL_23_896 ();
 FILLCELL_X32 FILLCELL_23_928 ();
 FILLCELL_X32 FILLCELL_23_960 ();
 FILLCELL_X32 FILLCELL_23_992 ();
 FILLCELL_X32 FILLCELL_23_1024 ();
 FILLCELL_X32 FILLCELL_23_1056 ();
 FILLCELL_X32 FILLCELL_23_1088 ();
 FILLCELL_X32 FILLCELL_23_1120 ();
 FILLCELL_X32 FILLCELL_23_1152 ();
 FILLCELL_X32 FILLCELL_23_1184 ();
 FILLCELL_X32 FILLCELL_23_1216 ();
 FILLCELL_X32 FILLCELL_23_1248 ();
 FILLCELL_X32 FILLCELL_23_1280 ();
 FILLCELL_X32 FILLCELL_23_1312 ();
 FILLCELL_X32 FILLCELL_23_1344 ();
 FILLCELL_X32 FILLCELL_23_1376 ();
 FILLCELL_X32 FILLCELL_23_1408 ();
 FILLCELL_X32 FILLCELL_23_1440 ();
 FILLCELL_X32 FILLCELL_23_1472 ();
 FILLCELL_X32 FILLCELL_23_1504 ();
 FILLCELL_X32 FILLCELL_23_1536 ();
 FILLCELL_X32 FILLCELL_23_1568 ();
 FILLCELL_X32 FILLCELL_23_1600 ();
 FILLCELL_X32 FILLCELL_23_1632 ();
 FILLCELL_X32 FILLCELL_23_1664 ();
 FILLCELL_X32 FILLCELL_23_1696 ();
 FILLCELL_X32 FILLCELL_23_1728 ();
 FILLCELL_X32 FILLCELL_23_1760 ();
 FILLCELL_X32 FILLCELL_23_1792 ();
 FILLCELL_X32 FILLCELL_23_1824 ();
 FILLCELL_X32 FILLCELL_23_1856 ();
 FILLCELL_X8 FILLCELL_23_1888 ();
 FILLCELL_X1 FILLCELL_23_1896 ();
 FILLCELL_X32 FILLCELL_24_0 ();
 FILLCELL_X32 FILLCELL_24_32 ();
 FILLCELL_X32 FILLCELL_24_64 ();
 FILLCELL_X32 FILLCELL_24_96 ();
 FILLCELL_X32 FILLCELL_24_128 ();
 FILLCELL_X32 FILLCELL_24_160 ();
 FILLCELL_X32 FILLCELL_24_192 ();
 FILLCELL_X32 FILLCELL_24_224 ();
 FILLCELL_X32 FILLCELL_24_256 ();
 FILLCELL_X32 FILLCELL_24_288 ();
 FILLCELL_X32 FILLCELL_24_320 ();
 FILLCELL_X32 FILLCELL_24_352 ();
 FILLCELL_X32 FILLCELL_24_384 ();
 FILLCELL_X32 FILLCELL_24_416 ();
 FILLCELL_X32 FILLCELL_24_448 ();
 FILLCELL_X32 FILLCELL_24_480 ();
 FILLCELL_X32 FILLCELL_24_512 ();
 FILLCELL_X32 FILLCELL_24_544 ();
 FILLCELL_X32 FILLCELL_24_576 ();
 FILLCELL_X32 FILLCELL_24_608 ();
 FILLCELL_X32 FILLCELL_24_640 ();
 FILLCELL_X32 FILLCELL_24_672 ();
 FILLCELL_X32 FILLCELL_24_704 ();
 FILLCELL_X32 FILLCELL_24_736 ();
 FILLCELL_X32 FILLCELL_24_768 ();
 FILLCELL_X32 FILLCELL_24_800 ();
 FILLCELL_X32 FILLCELL_24_832 ();
 FILLCELL_X32 FILLCELL_24_864 ();
 FILLCELL_X32 FILLCELL_24_896 ();
 FILLCELL_X32 FILLCELL_24_928 ();
 FILLCELL_X32 FILLCELL_24_960 ();
 FILLCELL_X32 FILLCELL_24_992 ();
 FILLCELL_X32 FILLCELL_24_1024 ();
 FILLCELL_X32 FILLCELL_24_1056 ();
 FILLCELL_X32 FILLCELL_24_1088 ();
 FILLCELL_X32 FILLCELL_24_1120 ();
 FILLCELL_X32 FILLCELL_24_1152 ();
 FILLCELL_X32 FILLCELL_24_1184 ();
 FILLCELL_X32 FILLCELL_24_1216 ();
 FILLCELL_X32 FILLCELL_24_1248 ();
 FILLCELL_X32 FILLCELL_24_1280 ();
 FILLCELL_X32 FILLCELL_24_1312 ();
 FILLCELL_X32 FILLCELL_24_1344 ();
 FILLCELL_X32 FILLCELL_24_1376 ();
 FILLCELL_X32 FILLCELL_24_1408 ();
 FILLCELL_X32 FILLCELL_24_1440 ();
 FILLCELL_X32 FILLCELL_24_1472 ();
 FILLCELL_X32 FILLCELL_24_1504 ();
 FILLCELL_X32 FILLCELL_24_1536 ();
 FILLCELL_X32 FILLCELL_24_1568 ();
 FILLCELL_X32 FILLCELL_24_1600 ();
 FILLCELL_X32 FILLCELL_24_1632 ();
 FILLCELL_X32 FILLCELL_24_1664 ();
 FILLCELL_X32 FILLCELL_24_1696 ();
 FILLCELL_X32 FILLCELL_24_1728 ();
 FILLCELL_X32 FILLCELL_24_1760 ();
 FILLCELL_X32 FILLCELL_24_1792 ();
 FILLCELL_X32 FILLCELL_24_1824 ();
 FILLCELL_X32 FILLCELL_24_1856 ();
 FILLCELL_X8 FILLCELL_24_1888 ();
 FILLCELL_X1 FILLCELL_24_1896 ();
 FILLCELL_X32 FILLCELL_25_0 ();
 FILLCELL_X32 FILLCELL_25_32 ();
 FILLCELL_X32 FILLCELL_25_64 ();
 FILLCELL_X32 FILLCELL_25_96 ();
 FILLCELL_X32 FILLCELL_25_128 ();
 FILLCELL_X32 FILLCELL_25_160 ();
 FILLCELL_X32 FILLCELL_25_192 ();
 FILLCELL_X32 FILLCELL_25_224 ();
 FILLCELL_X32 FILLCELL_25_256 ();
 FILLCELL_X32 FILLCELL_25_288 ();
 FILLCELL_X32 FILLCELL_25_320 ();
 FILLCELL_X32 FILLCELL_25_352 ();
 FILLCELL_X32 FILLCELL_25_384 ();
 FILLCELL_X32 FILLCELL_25_416 ();
 FILLCELL_X32 FILLCELL_25_448 ();
 FILLCELL_X32 FILLCELL_25_480 ();
 FILLCELL_X32 FILLCELL_25_512 ();
 FILLCELL_X32 FILLCELL_25_544 ();
 FILLCELL_X32 FILLCELL_25_576 ();
 FILLCELL_X32 FILLCELL_25_608 ();
 FILLCELL_X32 FILLCELL_25_640 ();
 FILLCELL_X32 FILLCELL_25_672 ();
 FILLCELL_X32 FILLCELL_25_704 ();
 FILLCELL_X32 FILLCELL_25_736 ();
 FILLCELL_X32 FILLCELL_25_768 ();
 FILLCELL_X32 FILLCELL_25_800 ();
 FILLCELL_X32 FILLCELL_25_832 ();
 FILLCELL_X32 FILLCELL_25_864 ();
 FILLCELL_X32 FILLCELL_25_896 ();
 FILLCELL_X32 FILLCELL_25_928 ();
 FILLCELL_X32 FILLCELL_25_960 ();
 FILLCELL_X32 FILLCELL_25_992 ();
 FILLCELL_X32 FILLCELL_25_1024 ();
 FILLCELL_X32 FILLCELL_25_1056 ();
 FILLCELL_X32 FILLCELL_25_1088 ();
 FILLCELL_X32 FILLCELL_25_1120 ();
 FILLCELL_X32 FILLCELL_25_1152 ();
 FILLCELL_X32 FILLCELL_25_1184 ();
 FILLCELL_X32 FILLCELL_25_1216 ();
 FILLCELL_X32 FILLCELL_25_1248 ();
 FILLCELL_X32 FILLCELL_25_1280 ();
 FILLCELL_X32 FILLCELL_25_1312 ();
 FILLCELL_X32 FILLCELL_25_1344 ();
 FILLCELL_X32 FILLCELL_25_1376 ();
 FILLCELL_X32 FILLCELL_25_1408 ();
 FILLCELL_X32 FILLCELL_25_1440 ();
 FILLCELL_X32 FILLCELL_25_1472 ();
 FILLCELL_X32 FILLCELL_25_1504 ();
 FILLCELL_X32 FILLCELL_25_1536 ();
 FILLCELL_X32 FILLCELL_25_1568 ();
 FILLCELL_X32 FILLCELL_25_1600 ();
 FILLCELL_X32 FILLCELL_25_1632 ();
 FILLCELL_X32 FILLCELL_25_1664 ();
 FILLCELL_X32 FILLCELL_25_1696 ();
 FILLCELL_X32 FILLCELL_25_1728 ();
 FILLCELL_X32 FILLCELL_25_1760 ();
 FILLCELL_X32 FILLCELL_25_1792 ();
 FILLCELL_X32 FILLCELL_25_1824 ();
 FILLCELL_X32 FILLCELL_25_1856 ();
 FILLCELL_X8 FILLCELL_25_1888 ();
 FILLCELL_X1 FILLCELL_25_1896 ();
 FILLCELL_X32 FILLCELL_26_0 ();
 FILLCELL_X32 FILLCELL_26_32 ();
 FILLCELL_X32 FILLCELL_26_64 ();
 FILLCELL_X32 FILLCELL_26_96 ();
 FILLCELL_X32 FILLCELL_26_128 ();
 FILLCELL_X32 FILLCELL_26_160 ();
 FILLCELL_X32 FILLCELL_26_192 ();
 FILLCELL_X32 FILLCELL_26_224 ();
 FILLCELL_X32 FILLCELL_26_256 ();
 FILLCELL_X32 FILLCELL_26_288 ();
 FILLCELL_X32 FILLCELL_26_320 ();
 FILLCELL_X32 FILLCELL_26_352 ();
 FILLCELL_X32 FILLCELL_26_384 ();
 FILLCELL_X32 FILLCELL_26_416 ();
 FILLCELL_X32 FILLCELL_26_448 ();
 FILLCELL_X32 FILLCELL_26_480 ();
 FILLCELL_X32 FILLCELL_26_512 ();
 FILLCELL_X32 FILLCELL_26_544 ();
 FILLCELL_X32 FILLCELL_26_576 ();
 FILLCELL_X32 FILLCELL_26_608 ();
 FILLCELL_X32 FILLCELL_26_640 ();
 FILLCELL_X32 FILLCELL_26_672 ();
 FILLCELL_X32 FILLCELL_26_704 ();
 FILLCELL_X32 FILLCELL_26_736 ();
 FILLCELL_X32 FILLCELL_26_768 ();
 FILLCELL_X32 FILLCELL_26_800 ();
 FILLCELL_X32 FILLCELL_26_832 ();
 FILLCELL_X32 FILLCELL_26_864 ();
 FILLCELL_X32 FILLCELL_26_896 ();
 FILLCELL_X32 FILLCELL_26_928 ();
 FILLCELL_X32 FILLCELL_26_960 ();
 FILLCELL_X32 FILLCELL_26_992 ();
 FILLCELL_X32 FILLCELL_26_1024 ();
 FILLCELL_X32 FILLCELL_26_1056 ();
 FILLCELL_X32 FILLCELL_26_1088 ();
 FILLCELL_X32 FILLCELL_26_1120 ();
 FILLCELL_X32 FILLCELL_26_1152 ();
 FILLCELL_X32 FILLCELL_26_1184 ();
 FILLCELL_X32 FILLCELL_26_1216 ();
 FILLCELL_X32 FILLCELL_26_1248 ();
 FILLCELL_X32 FILLCELL_26_1280 ();
 FILLCELL_X32 FILLCELL_26_1312 ();
 FILLCELL_X32 FILLCELL_26_1344 ();
 FILLCELL_X32 FILLCELL_26_1376 ();
 FILLCELL_X32 FILLCELL_26_1408 ();
 FILLCELL_X32 FILLCELL_26_1440 ();
 FILLCELL_X32 FILLCELL_26_1472 ();
 FILLCELL_X32 FILLCELL_26_1504 ();
 FILLCELL_X32 FILLCELL_26_1536 ();
 FILLCELL_X32 FILLCELL_26_1568 ();
 FILLCELL_X32 FILLCELL_26_1600 ();
 FILLCELL_X32 FILLCELL_26_1632 ();
 FILLCELL_X32 FILLCELL_26_1664 ();
 FILLCELL_X32 FILLCELL_26_1696 ();
 FILLCELL_X32 FILLCELL_26_1728 ();
 FILLCELL_X32 FILLCELL_26_1760 ();
 FILLCELL_X32 FILLCELL_26_1792 ();
 FILLCELL_X32 FILLCELL_26_1824 ();
 FILLCELL_X32 FILLCELL_26_1856 ();
 FILLCELL_X8 FILLCELL_26_1888 ();
 FILLCELL_X1 FILLCELL_26_1896 ();
 FILLCELL_X32 FILLCELL_27_0 ();
 FILLCELL_X32 FILLCELL_27_32 ();
 FILLCELL_X32 FILLCELL_27_64 ();
 FILLCELL_X32 FILLCELL_27_96 ();
 FILLCELL_X32 FILLCELL_27_128 ();
 FILLCELL_X32 FILLCELL_27_160 ();
 FILLCELL_X32 FILLCELL_27_192 ();
 FILLCELL_X32 FILLCELL_27_224 ();
 FILLCELL_X32 FILLCELL_27_256 ();
 FILLCELL_X32 FILLCELL_27_288 ();
 FILLCELL_X32 FILLCELL_27_320 ();
 FILLCELL_X32 FILLCELL_27_352 ();
 FILLCELL_X32 FILLCELL_27_384 ();
 FILLCELL_X32 FILLCELL_27_416 ();
 FILLCELL_X32 FILLCELL_27_448 ();
 FILLCELL_X32 FILLCELL_27_480 ();
 FILLCELL_X32 FILLCELL_27_512 ();
 FILLCELL_X32 FILLCELL_27_544 ();
 FILLCELL_X32 FILLCELL_27_576 ();
 FILLCELL_X32 FILLCELL_27_608 ();
 FILLCELL_X32 FILLCELL_27_640 ();
 FILLCELL_X32 FILLCELL_27_672 ();
 FILLCELL_X32 FILLCELL_27_704 ();
 FILLCELL_X32 FILLCELL_27_736 ();
 FILLCELL_X32 FILLCELL_27_768 ();
 FILLCELL_X32 FILLCELL_27_800 ();
 FILLCELL_X32 FILLCELL_27_832 ();
 FILLCELL_X32 FILLCELL_27_864 ();
 FILLCELL_X32 FILLCELL_27_896 ();
 FILLCELL_X32 FILLCELL_27_928 ();
 FILLCELL_X32 FILLCELL_27_960 ();
 FILLCELL_X32 FILLCELL_27_992 ();
 FILLCELL_X32 FILLCELL_27_1024 ();
 FILLCELL_X32 FILLCELL_27_1056 ();
 FILLCELL_X32 FILLCELL_27_1088 ();
 FILLCELL_X32 FILLCELL_27_1120 ();
 FILLCELL_X32 FILLCELL_27_1152 ();
 FILLCELL_X32 FILLCELL_27_1184 ();
 FILLCELL_X32 FILLCELL_27_1216 ();
 FILLCELL_X32 FILLCELL_27_1248 ();
 FILLCELL_X32 FILLCELL_27_1280 ();
 FILLCELL_X32 FILLCELL_27_1312 ();
 FILLCELL_X32 FILLCELL_27_1344 ();
 FILLCELL_X32 FILLCELL_27_1376 ();
 FILLCELL_X32 FILLCELL_27_1408 ();
 FILLCELL_X32 FILLCELL_27_1440 ();
 FILLCELL_X32 FILLCELL_27_1472 ();
 FILLCELL_X32 FILLCELL_27_1504 ();
 FILLCELL_X32 FILLCELL_27_1536 ();
 FILLCELL_X32 FILLCELL_27_1568 ();
 FILLCELL_X32 FILLCELL_27_1600 ();
 FILLCELL_X32 FILLCELL_27_1632 ();
 FILLCELL_X32 FILLCELL_27_1664 ();
 FILLCELL_X32 FILLCELL_27_1696 ();
 FILLCELL_X32 FILLCELL_27_1728 ();
 FILLCELL_X32 FILLCELL_27_1760 ();
 FILLCELL_X32 FILLCELL_27_1792 ();
 FILLCELL_X32 FILLCELL_27_1824 ();
 FILLCELL_X32 FILLCELL_27_1856 ();
 FILLCELL_X8 FILLCELL_27_1888 ();
 FILLCELL_X1 FILLCELL_27_1896 ();
 FILLCELL_X32 FILLCELL_28_0 ();
 FILLCELL_X32 FILLCELL_28_32 ();
 FILLCELL_X32 FILLCELL_28_64 ();
 FILLCELL_X32 FILLCELL_28_96 ();
 FILLCELL_X32 FILLCELL_28_128 ();
 FILLCELL_X32 FILLCELL_28_160 ();
 FILLCELL_X32 FILLCELL_28_192 ();
 FILLCELL_X32 FILLCELL_28_224 ();
 FILLCELL_X32 FILLCELL_28_256 ();
 FILLCELL_X32 FILLCELL_28_288 ();
 FILLCELL_X32 FILLCELL_28_320 ();
 FILLCELL_X32 FILLCELL_28_352 ();
 FILLCELL_X32 FILLCELL_28_384 ();
 FILLCELL_X32 FILLCELL_28_416 ();
 FILLCELL_X32 FILLCELL_28_448 ();
 FILLCELL_X32 FILLCELL_28_480 ();
 FILLCELL_X32 FILLCELL_28_512 ();
 FILLCELL_X32 FILLCELL_28_544 ();
 FILLCELL_X32 FILLCELL_28_576 ();
 FILLCELL_X32 FILLCELL_28_608 ();
 FILLCELL_X32 FILLCELL_28_640 ();
 FILLCELL_X32 FILLCELL_28_672 ();
 FILLCELL_X32 FILLCELL_28_704 ();
 FILLCELL_X32 FILLCELL_28_736 ();
 FILLCELL_X32 FILLCELL_28_768 ();
 FILLCELL_X32 FILLCELL_28_800 ();
 FILLCELL_X32 FILLCELL_28_832 ();
 FILLCELL_X32 FILLCELL_28_864 ();
 FILLCELL_X32 FILLCELL_28_896 ();
 FILLCELL_X32 FILLCELL_28_928 ();
 FILLCELL_X32 FILLCELL_28_960 ();
 FILLCELL_X32 FILLCELL_28_992 ();
 FILLCELL_X32 FILLCELL_28_1024 ();
 FILLCELL_X32 FILLCELL_28_1056 ();
 FILLCELL_X32 FILLCELL_28_1088 ();
 FILLCELL_X32 FILLCELL_28_1120 ();
 FILLCELL_X32 FILLCELL_28_1152 ();
 FILLCELL_X32 FILLCELL_28_1184 ();
 FILLCELL_X32 FILLCELL_28_1216 ();
 FILLCELL_X32 FILLCELL_28_1248 ();
 FILLCELL_X32 FILLCELL_28_1280 ();
 FILLCELL_X32 FILLCELL_28_1312 ();
 FILLCELL_X32 FILLCELL_28_1344 ();
 FILLCELL_X32 FILLCELL_28_1376 ();
 FILLCELL_X32 FILLCELL_28_1408 ();
 FILLCELL_X32 FILLCELL_28_1440 ();
 FILLCELL_X32 FILLCELL_28_1472 ();
 FILLCELL_X32 FILLCELL_28_1504 ();
 FILLCELL_X32 FILLCELL_28_1536 ();
 FILLCELL_X32 FILLCELL_28_1568 ();
 FILLCELL_X32 FILLCELL_28_1600 ();
 FILLCELL_X32 FILLCELL_28_1632 ();
 FILLCELL_X32 FILLCELL_28_1664 ();
 FILLCELL_X32 FILLCELL_28_1696 ();
 FILLCELL_X32 FILLCELL_28_1728 ();
 FILLCELL_X32 FILLCELL_28_1760 ();
 FILLCELL_X32 FILLCELL_28_1792 ();
 FILLCELL_X32 FILLCELL_28_1824 ();
 FILLCELL_X32 FILLCELL_28_1856 ();
 FILLCELL_X8 FILLCELL_28_1888 ();
 FILLCELL_X1 FILLCELL_28_1896 ();
 FILLCELL_X32 FILLCELL_29_0 ();
 FILLCELL_X32 FILLCELL_29_32 ();
 FILLCELL_X32 FILLCELL_29_64 ();
 FILLCELL_X32 FILLCELL_29_96 ();
 FILLCELL_X32 FILLCELL_29_128 ();
 FILLCELL_X32 FILLCELL_29_160 ();
 FILLCELL_X32 FILLCELL_29_192 ();
 FILLCELL_X32 FILLCELL_29_224 ();
 FILLCELL_X32 FILLCELL_29_256 ();
 FILLCELL_X32 FILLCELL_29_288 ();
 FILLCELL_X32 FILLCELL_29_320 ();
 FILLCELL_X32 FILLCELL_29_352 ();
 FILLCELL_X32 FILLCELL_29_384 ();
 FILLCELL_X32 FILLCELL_29_416 ();
 FILLCELL_X32 FILLCELL_29_448 ();
 FILLCELL_X32 FILLCELL_29_480 ();
 FILLCELL_X32 FILLCELL_29_512 ();
 FILLCELL_X32 FILLCELL_29_544 ();
 FILLCELL_X32 FILLCELL_29_576 ();
 FILLCELL_X32 FILLCELL_29_608 ();
 FILLCELL_X32 FILLCELL_29_640 ();
 FILLCELL_X32 FILLCELL_29_672 ();
 FILLCELL_X32 FILLCELL_29_704 ();
 FILLCELL_X32 FILLCELL_29_736 ();
 FILLCELL_X32 FILLCELL_29_768 ();
 FILLCELL_X32 FILLCELL_29_800 ();
 FILLCELL_X32 FILLCELL_29_832 ();
 FILLCELL_X32 FILLCELL_29_864 ();
 FILLCELL_X32 FILLCELL_29_896 ();
 FILLCELL_X32 FILLCELL_29_928 ();
 FILLCELL_X32 FILLCELL_29_960 ();
 FILLCELL_X32 FILLCELL_29_992 ();
 FILLCELL_X32 FILLCELL_29_1024 ();
 FILLCELL_X32 FILLCELL_29_1056 ();
 FILLCELL_X32 FILLCELL_29_1088 ();
 FILLCELL_X32 FILLCELL_29_1120 ();
 FILLCELL_X32 FILLCELL_29_1152 ();
 FILLCELL_X32 FILLCELL_29_1184 ();
 FILLCELL_X32 FILLCELL_29_1216 ();
 FILLCELL_X32 FILLCELL_29_1248 ();
 FILLCELL_X32 FILLCELL_29_1280 ();
 FILLCELL_X32 FILLCELL_29_1312 ();
 FILLCELL_X32 FILLCELL_29_1344 ();
 FILLCELL_X32 FILLCELL_29_1376 ();
 FILLCELL_X32 FILLCELL_29_1408 ();
 FILLCELL_X32 FILLCELL_29_1440 ();
 FILLCELL_X32 FILLCELL_29_1472 ();
 FILLCELL_X32 FILLCELL_29_1504 ();
 FILLCELL_X32 FILLCELL_29_1536 ();
 FILLCELL_X32 FILLCELL_29_1568 ();
 FILLCELL_X32 FILLCELL_29_1600 ();
 FILLCELL_X32 FILLCELL_29_1632 ();
 FILLCELL_X32 FILLCELL_29_1664 ();
 FILLCELL_X32 FILLCELL_29_1696 ();
 FILLCELL_X32 FILLCELL_29_1728 ();
 FILLCELL_X32 FILLCELL_29_1760 ();
 FILLCELL_X32 FILLCELL_29_1792 ();
 FILLCELL_X32 FILLCELL_29_1824 ();
 FILLCELL_X32 FILLCELL_29_1856 ();
 FILLCELL_X8 FILLCELL_29_1888 ();
 FILLCELL_X1 FILLCELL_29_1896 ();
 FILLCELL_X32 FILLCELL_30_0 ();
 FILLCELL_X32 FILLCELL_30_32 ();
 FILLCELL_X32 FILLCELL_30_64 ();
 FILLCELL_X32 FILLCELL_30_96 ();
 FILLCELL_X32 FILLCELL_30_128 ();
 FILLCELL_X32 FILLCELL_30_160 ();
 FILLCELL_X32 FILLCELL_30_192 ();
 FILLCELL_X32 FILLCELL_30_224 ();
 FILLCELL_X32 FILLCELL_30_256 ();
 FILLCELL_X32 FILLCELL_30_288 ();
 FILLCELL_X32 FILLCELL_30_320 ();
 FILLCELL_X32 FILLCELL_30_352 ();
 FILLCELL_X32 FILLCELL_30_384 ();
 FILLCELL_X32 FILLCELL_30_416 ();
 FILLCELL_X32 FILLCELL_30_448 ();
 FILLCELL_X32 FILLCELL_30_480 ();
 FILLCELL_X32 FILLCELL_30_512 ();
 FILLCELL_X32 FILLCELL_30_544 ();
 FILLCELL_X32 FILLCELL_30_576 ();
 FILLCELL_X32 FILLCELL_30_608 ();
 FILLCELL_X32 FILLCELL_30_640 ();
 FILLCELL_X32 FILLCELL_30_672 ();
 FILLCELL_X32 FILLCELL_30_704 ();
 FILLCELL_X32 FILLCELL_30_736 ();
 FILLCELL_X32 FILLCELL_30_768 ();
 FILLCELL_X32 FILLCELL_30_800 ();
 FILLCELL_X32 FILLCELL_30_832 ();
 FILLCELL_X32 FILLCELL_30_864 ();
 FILLCELL_X32 FILLCELL_30_896 ();
 FILLCELL_X32 FILLCELL_30_928 ();
 FILLCELL_X32 FILLCELL_30_960 ();
 FILLCELL_X32 FILLCELL_30_992 ();
 FILLCELL_X32 FILLCELL_30_1024 ();
 FILLCELL_X32 FILLCELL_30_1056 ();
 FILLCELL_X32 FILLCELL_30_1088 ();
 FILLCELL_X32 FILLCELL_30_1120 ();
 FILLCELL_X32 FILLCELL_30_1152 ();
 FILLCELL_X32 FILLCELL_30_1184 ();
 FILLCELL_X32 FILLCELL_30_1216 ();
 FILLCELL_X32 FILLCELL_30_1248 ();
 FILLCELL_X32 FILLCELL_30_1280 ();
 FILLCELL_X32 FILLCELL_30_1312 ();
 FILLCELL_X32 FILLCELL_30_1344 ();
 FILLCELL_X32 FILLCELL_30_1376 ();
 FILLCELL_X32 FILLCELL_30_1408 ();
 FILLCELL_X32 FILLCELL_30_1440 ();
 FILLCELL_X32 FILLCELL_30_1472 ();
 FILLCELL_X32 FILLCELL_30_1504 ();
 FILLCELL_X32 FILLCELL_30_1536 ();
 FILLCELL_X32 FILLCELL_30_1568 ();
 FILLCELL_X32 FILLCELL_30_1600 ();
 FILLCELL_X32 FILLCELL_30_1632 ();
 FILLCELL_X32 FILLCELL_30_1664 ();
 FILLCELL_X32 FILLCELL_30_1696 ();
 FILLCELL_X32 FILLCELL_30_1728 ();
 FILLCELL_X32 FILLCELL_30_1760 ();
 FILLCELL_X32 FILLCELL_30_1792 ();
 FILLCELL_X32 FILLCELL_30_1824 ();
 FILLCELL_X32 FILLCELL_30_1856 ();
 FILLCELL_X8 FILLCELL_30_1888 ();
 FILLCELL_X1 FILLCELL_30_1896 ();
 FILLCELL_X32 FILLCELL_31_0 ();
 FILLCELL_X32 FILLCELL_31_32 ();
 FILLCELL_X32 FILLCELL_31_64 ();
 FILLCELL_X32 FILLCELL_31_96 ();
 FILLCELL_X32 FILLCELL_31_128 ();
 FILLCELL_X32 FILLCELL_31_160 ();
 FILLCELL_X32 FILLCELL_31_192 ();
 FILLCELL_X32 FILLCELL_31_224 ();
 FILLCELL_X32 FILLCELL_31_256 ();
 FILLCELL_X32 FILLCELL_31_288 ();
 FILLCELL_X32 FILLCELL_31_320 ();
 FILLCELL_X32 FILLCELL_31_352 ();
 FILLCELL_X32 FILLCELL_31_384 ();
 FILLCELL_X32 FILLCELL_31_416 ();
 FILLCELL_X32 FILLCELL_31_448 ();
 FILLCELL_X32 FILLCELL_31_480 ();
 FILLCELL_X32 FILLCELL_31_512 ();
 FILLCELL_X32 FILLCELL_31_544 ();
 FILLCELL_X32 FILLCELL_31_576 ();
 FILLCELL_X32 FILLCELL_31_608 ();
 FILLCELL_X32 FILLCELL_31_640 ();
 FILLCELL_X32 FILLCELL_31_672 ();
 FILLCELL_X32 FILLCELL_31_704 ();
 FILLCELL_X32 FILLCELL_31_736 ();
 FILLCELL_X32 FILLCELL_31_768 ();
 FILLCELL_X32 FILLCELL_31_800 ();
 FILLCELL_X32 FILLCELL_31_832 ();
 FILLCELL_X32 FILLCELL_31_864 ();
 FILLCELL_X32 FILLCELL_31_896 ();
 FILLCELL_X32 FILLCELL_31_928 ();
 FILLCELL_X32 FILLCELL_31_960 ();
 FILLCELL_X32 FILLCELL_31_992 ();
 FILLCELL_X32 FILLCELL_31_1024 ();
 FILLCELL_X32 FILLCELL_31_1056 ();
 FILLCELL_X32 FILLCELL_31_1088 ();
 FILLCELL_X32 FILLCELL_31_1120 ();
 FILLCELL_X32 FILLCELL_31_1152 ();
 FILLCELL_X32 FILLCELL_31_1184 ();
 FILLCELL_X32 FILLCELL_31_1216 ();
 FILLCELL_X32 FILLCELL_31_1248 ();
 FILLCELL_X32 FILLCELL_31_1280 ();
 FILLCELL_X32 FILLCELL_31_1312 ();
 FILLCELL_X32 FILLCELL_31_1344 ();
 FILLCELL_X32 FILLCELL_31_1376 ();
 FILLCELL_X32 FILLCELL_31_1408 ();
 FILLCELL_X32 FILLCELL_31_1440 ();
 FILLCELL_X32 FILLCELL_31_1472 ();
 FILLCELL_X32 FILLCELL_31_1504 ();
 FILLCELL_X32 FILLCELL_31_1536 ();
 FILLCELL_X32 FILLCELL_31_1568 ();
 FILLCELL_X32 FILLCELL_31_1600 ();
 FILLCELL_X32 FILLCELL_31_1632 ();
 FILLCELL_X32 FILLCELL_31_1664 ();
 FILLCELL_X32 FILLCELL_31_1696 ();
 FILLCELL_X32 FILLCELL_31_1728 ();
 FILLCELL_X32 FILLCELL_31_1760 ();
 FILLCELL_X32 FILLCELL_31_1792 ();
 FILLCELL_X32 FILLCELL_31_1824 ();
 FILLCELL_X32 FILLCELL_31_1856 ();
 FILLCELL_X8 FILLCELL_31_1888 ();
 FILLCELL_X1 FILLCELL_31_1896 ();
 FILLCELL_X32 FILLCELL_32_0 ();
 FILLCELL_X32 FILLCELL_32_32 ();
 FILLCELL_X32 FILLCELL_32_64 ();
 FILLCELL_X32 FILLCELL_32_96 ();
 FILLCELL_X32 FILLCELL_32_128 ();
 FILLCELL_X32 FILLCELL_32_160 ();
 FILLCELL_X32 FILLCELL_32_192 ();
 FILLCELL_X32 FILLCELL_32_224 ();
 FILLCELL_X32 FILLCELL_32_256 ();
 FILLCELL_X32 FILLCELL_32_288 ();
 FILLCELL_X32 FILLCELL_32_320 ();
 FILLCELL_X32 FILLCELL_32_352 ();
 FILLCELL_X32 FILLCELL_32_384 ();
 FILLCELL_X32 FILLCELL_32_416 ();
 FILLCELL_X32 FILLCELL_32_448 ();
 FILLCELL_X32 FILLCELL_32_480 ();
 FILLCELL_X32 FILLCELL_32_512 ();
 FILLCELL_X32 FILLCELL_32_544 ();
 FILLCELL_X32 FILLCELL_32_576 ();
 FILLCELL_X32 FILLCELL_32_608 ();
 FILLCELL_X32 FILLCELL_32_640 ();
 FILLCELL_X32 FILLCELL_32_672 ();
 FILLCELL_X32 FILLCELL_32_704 ();
 FILLCELL_X32 FILLCELL_32_736 ();
 FILLCELL_X32 FILLCELL_32_768 ();
 FILLCELL_X32 FILLCELL_32_800 ();
 FILLCELL_X32 FILLCELL_32_832 ();
 FILLCELL_X32 FILLCELL_32_864 ();
 FILLCELL_X32 FILLCELL_32_896 ();
 FILLCELL_X32 FILLCELL_32_928 ();
 FILLCELL_X32 FILLCELL_32_960 ();
 FILLCELL_X32 FILLCELL_32_992 ();
 FILLCELL_X32 FILLCELL_32_1024 ();
 FILLCELL_X32 FILLCELL_32_1056 ();
 FILLCELL_X32 FILLCELL_32_1088 ();
 FILLCELL_X32 FILLCELL_32_1120 ();
 FILLCELL_X32 FILLCELL_32_1152 ();
 FILLCELL_X32 FILLCELL_32_1184 ();
 FILLCELL_X32 FILLCELL_32_1216 ();
 FILLCELL_X32 FILLCELL_32_1248 ();
 FILLCELL_X32 FILLCELL_32_1280 ();
 FILLCELL_X32 FILLCELL_32_1312 ();
 FILLCELL_X32 FILLCELL_32_1344 ();
 FILLCELL_X32 FILLCELL_32_1376 ();
 FILLCELL_X32 FILLCELL_32_1408 ();
 FILLCELL_X32 FILLCELL_32_1440 ();
 FILLCELL_X32 FILLCELL_32_1472 ();
 FILLCELL_X32 FILLCELL_32_1504 ();
 FILLCELL_X32 FILLCELL_32_1536 ();
 FILLCELL_X32 FILLCELL_32_1568 ();
 FILLCELL_X32 FILLCELL_32_1600 ();
 FILLCELL_X32 FILLCELL_32_1632 ();
 FILLCELL_X32 FILLCELL_32_1664 ();
 FILLCELL_X32 FILLCELL_32_1696 ();
 FILLCELL_X32 FILLCELL_32_1728 ();
 FILLCELL_X32 FILLCELL_32_1760 ();
 FILLCELL_X32 FILLCELL_32_1792 ();
 FILLCELL_X32 FILLCELL_32_1824 ();
 FILLCELL_X32 FILLCELL_32_1856 ();
 FILLCELL_X8 FILLCELL_32_1888 ();
 FILLCELL_X1 FILLCELL_32_1896 ();
 FILLCELL_X32 FILLCELL_33_0 ();
 FILLCELL_X32 FILLCELL_33_32 ();
 FILLCELL_X32 FILLCELL_33_64 ();
 FILLCELL_X32 FILLCELL_33_96 ();
 FILLCELL_X32 FILLCELL_33_128 ();
 FILLCELL_X32 FILLCELL_33_160 ();
 FILLCELL_X32 FILLCELL_33_192 ();
 FILLCELL_X32 FILLCELL_33_224 ();
 FILLCELL_X32 FILLCELL_33_256 ();
 FILLCELL_X32 FILLCELL_33_288 ();
 FILLCELL_X32 FILLCELL_33_320 ();
 FILLCELL_X32 FILLCELL_33_352 ();
 FILLCELL_X32 FILLCELL_33_384 ();
 FILLCELL_X32 FILLCELL_33_416 ();
 FILLCELL_X32 FILLCELL_33_448 ();
 FILLCELL_X32 FILLCELL_33_480 ();
 FILLCELL_X32 FILLCELL_33_512 ();
 FILLCELL_X32 FILLCELL_33_544 ();
 FILLCELL_X32 FILLCELL_33_576 ();
 FILLCELL_X32 FILLCELL_33_608 ();
 FILLCELL_X32 FILLCELL_33_640 ();
 FILLCELL_X32 FILLCELL_33_672 ();
 FILLCELL_X32 FILLCELL_33_704 ();
 FILLCELL_X32 FILLCELL_33_736 ();
 FILLCELL_X32 FILLCELL_33_768 ();
 FILLCELL_X32 FILLCELL_33_800 ();
 FILLCELL_X32 FILLCELL_33_832 ();
 FILLCELL_X32 FILLCELL_33_864 ();
 FILLCELL_X32 FILLCELL_33_896 ();
 FILLCELL_X32 FILLCELL_33_928 ();
 FILLCELL_X32 FILLCELL_33_960 ();
 FILLCELL_X32 FILLCELL_33_992 ();
 FILLCELL_X32 FILLCELL_33_1024 ();
 FILLCELL_X32 FILLCELL_33_1056 ();
 FILLCELL_X32 FILLCELL_33_1088 ();
 FILLCELL_X32 FILLCELL_33_1120 ();
 FILLCELL_X32 FILLCELL_33_1152 ();
 FILLCELL_X32 FILLCELL_33_1184 ();
 FILLCELL_X32 FILLCELL_33_1216 ();
 FILLCELL_X32 FILLCELL_33_1248 ();
 FILLCELL_X32 FILLCELL_33_1280 ();
 FILLCELL_X32 FILLCELL_33_1312 ();
 FILLCELL_X32 FILLCELL_33_1344 ();
 FILLCELL_X32 FILLCELL_33_1376 ();
 FILLCELL_X32 FILLCELL_33_1408 ();
 FILLCELL_X32 FILLCELL_33_1440 ();
 FILLCELL_X32 FILLCELL_33_1472 ();
 FILLCELL_X32 FILLCELL_33_1504 ();
 FILLCELL_X32 FILLCELL_33_1536 ();
 FILLCELL_X32 FILLCELL_33_1568 ();
 FILLCELL_X32 FILLCELL_33_1600 ();
 FILLCELL_X32 FILLCELL_33_1632 ();
 FILLCELL_X32 FILLCELL_33_1664 ();
 FILLCELL_X32 FILLCELL_33_1696 ();
 FILLCELL_X32 FILLCELL_33_1728 ();
 FILLCELL_X32 FILLCELL_33_1760 ();
 FILLCELL_X32 FILLCELL_33_1792 ();
 FILLCELL_X32 FILLCELL_33_1824 ();
 FILLCELL_X32 FILLCELL_33_1856 ();
 FILLCELL_X8 FILLCELL_33_1888 ();
 FILLCELL_X1 FILLCELL_33_1896 ();
 FILLCELL_X32 FILLCELL_34_0 ();
 FILLCELL_X32 FILLCELL_34_32 ();
 FILLCELL_X32 FILLCELL_34_64 ();
 FILLCELL_X32 FILLCELL_34_96 ();
 FILLCELL_X32 FILLCELL_34_128 ();
 FILLCELL_X32 FILLCELL_34_160 ();
 FILLCELL_X32 FILLCELL_34_192 ();
 FILLCELL_X32 FILLCELL_34_224 ();
 FILLCELL_X32 FILLCELL_34_256 ();
 FILLCELL_X32 FILLCELL_34_288 ();
 FILLCELL_X32 FILLCELL_34_320 ();
 FILLCELL_X32 FILLCELL_34_352 ();
 FILLCELL_X32 FILLCELL_34_384 ();
 FILLCELL_X32 FILLCELL_34_416 ();
 FILLCELL_X32 FILLCELL_34_448 ();
 FILLCELL_X32 FILLCELL_34_480 ();
 FILLCELL_X32 FILLCELL_34_512 ();
 FILLCELL_X32 FILLCELL_34_544 ();
 FILLCELL_X32 FILLCELL_34_576 ();
 FILLCELL_X32 FILLCELL_34_608 ();
 FILLCELL_X32 FILLCELL_34_640 ();
 FILLCELL_X32 FILLCELL_34_672 ();
 FILLCELL_X32 FILLCELL_34_704 ();
 FILLCELL_X32 FILLCELL_34_736 ();
 FILLCELL_X32 FILLCELL_34_768 ();
 FILLCELL_X32 FILLCELL_34_800 ();
 FILLCELL_X32 FILLCELL_34_832 ();
 FILLCELL_X32 FILLCELL_34_864 ();
 FILLCELL_X32 FILLCELL_34_896 ();
 FILLCELL_X32 FILLCELL_34_928 ();
 FILLCELL_X32 FILLCELL_34_960 ();
 FILLCELL_X32 FILLCELL_34_992 ();
 FILLCELL_X32 FILLCELL_34_1024 ();
 FILLCELL_X32 FILLCELL_34_1056 ();
 FILLCELL_X32 FILLCELL_34_1088 ();
 FILLCELL_X32 FILLCELL_34_1120 ();
 FILLCELL_X32 FILLCELL_34_1152 ();
 FILLCELL_X32 FILLCELL_34_1184 ();
 FILLCELL_X32 FILLCELL_34_1216 ();
 FILLCELL_X32 FILLCELL_34_1248 ();
 FILLCELL_X32 FILLCELL_34_1280 ();
 FILLCELL_X32 FILLCELL_34_1312 ();
 FILLCELL_X32 FILLCELL_34_1344 ();
 FILLCELL_X32 FILLCELL_34_1376 ();
 FILLCELL_X32 FILLCELL_34_1408 ();
 FILLCELL_X32 FILLCELL_34_1440 ();
 FILLCELL_X32 FILLCELL_34_1472 ();
 FILLCELL_X32 FILLCELL_34_1504 ();
 FILLCELL_X32 FILLCELL_34_1536 ();
 FILLCELL_X32 FILLCELL_34_1568 ();
 FILLCELL_X32 FILLCELL_34_1600 ();
 FILLCELL_X32 FILLCELL_34_1632 ();
 FILLCELL_X32 FILLCELL_34_1664 ();
 FILLCELL_X32 FILLCELL_34_1696 ();
 FILLCELL_X32 FILLCELL_34_1728 ();
 FILLCELL_X32 FILLCELL_34_1760 ();
 FILLCELL_X32 FILLCELL_34_1792 ();
 FILLCELL_X32 FILLCELL_34_1824 ();
 FILLCELL_X32 FILLCELL_34_1856 ();
 FILLCELL_X8 FILLCELL_34_1888 ();
 FILLCELL_X1 FILLCELL_34_1896 ();
 FILLCELL_X32 FILLCELL_35_0 ();
 FILLCELL_X32 FILLCELL_35_32 ();
 FILLCELL_X32 FILLCELL_35_64 ();
 FILLCELL_X32 FILLCELL_35_96 ();
 FILLCELL_X32 FILLCELL_35_128 ();
 FILLCELL_X32 FILLCELL_35_160 ();
 FILLCELL_X32 FILLCELL_35_192 ();
 FILLCELL_X32 FILLCELL_35_224 ();
 FILLCELL_X32 FILLCELL_35_256 ();
 FILLCELL_X32 FILLCELL_35_288 ();
 FILLCELL_X32 FILLCELL_35_320 ();
 FILLCELL_X32 FILLCELL_35_352 ();
 FILLCELL_X32 FILLCELL_35_384 ();
 FILLCELL_X32 FILLCELL_35_416 ();
 FILLCELL_X32 FILLCELL_35_448 ();
 FILLCELL_X32 FILLCELL_35_480 ();
 FILLCELL_X32 FILLCELL_35_512 ();
 FILLCELL_X32 FILLCELL_35_544 ();
 FILLCELL_X32 FILLCELL_35_576 ();
 FILLCELL_X32 FILLCELL_35_608 ();
 FILLCELL_X32 FILLCELL_35_640 ();
 FILLCELL_X32 FILLCELL_35_672 ();
 FILLCELL_X32 FILLCELL_35_704 ();
 FILLCELL_X32 FILLCELL_35_736 ();
 FILLCELL_X32 FILLCELL_35_768 ();
 FILLCELL_X32 FILLCELL_35_800 ();
 FILLCELL_X32 FILLCELL_35_832 ();
 FILLCELL_X32 FILLCELL_35_864 ();
 FILLCELL_X32 FILLCELL_35_896 ();
 FILLCELL_X32 FILLCELL_35_928 ();
 FILLCELL_X32 FILLCELL_35_960 ();
 FILLCELL_X32 FILLCELL_35_992 ();
 FILLCELL_X32 FILLCELL_35_1024 ();
 FILLCELL_X32 FILLCELL_35_1056 ();
 FILLCELL_X32 FILLCELL_35_1088 ();
 FILLCELL_X32 FILLCELL_35_1120 ();
 FILLCELL_X32 FILLCELL_35_1152 ();
 FILLCELL_X32 FILLCELL_35_1184 ();
 FILLCELL_X32 FILLCELL_35_1216 ();
 FILLCELL_X32 FILLCELL_35_1248 ();
 FILLCELL_X32 FILLCELL_35_1280 ();
 FILLCELL_X32 FILLCELL_35_1312 ();
 FILLCELL_X32 FILLCELL_35_1344 ();
 FILLCELL_X32 FILLCELL_35_1376 ();
 FILLCELL_X32 FILLCELL_35_1408 ();
 FILLCELL_X32 FILLCELL_35_1440 ();
 FILLCELL_X32 FILLCELL_35_1472 ();
 FILLCELL_X32 FILLCELL_35_1504 ();
 FILLCELL_X32 FILLCELL_35_1536 ();
 FILLCELL_X32 FILLCELL_35_1568 ();
 FILLCELL_X32 FILLCELL_35_1600 ();
 FILLCELL_X32 FILLCELL_35_1632 ();
 FILLCELL_X32 FILLCELL_35_1664 ();
 FILLCELL_X32 FILLCELL_35_1696 ();
 FILLCELL_X32 FILLCELL_35_1728 ();
 FILLCELL_X32 FILLCELL_35_1760 ();
 FILLCELL_X32 FILLCELL_35_1792 ();
 FILLCELL_X32 FILLCELL_35_1824 ();
 FILLCELL_X32 FILLCELL_35_1856 ();
 FILLCELL_X8 FILLCELL_35_1888 ();
 FILLCELL_X1 FILLCELL_35_1896 ();
 FILLCELL_X32 FILLCELL_36_0 ();
 FILLCELL_X32 FILLCELL_36_32 ();
 FILLCELL_X32 FILLCELL_36_64 ();
 FILLCELL_X32 FILLCELL_36_96 ();
 FILLCELL_X32 FILLCELL_36_128 ();
 FILLCELL_X32 FILLCELL_36_160 ();
 FILLCELL_X32 FILLCELL_36_192 ();
 FILLCELL_X32 FILLCELL_36_224 ();
 FILLCELL_X32 FILLCELL_36_256 ();
 FILLCELL_X32 FILLCELL_36_288 ();
 FILLCELL_X32 FILLCELL_36_320 ();
 FILLCELL_X32 FILLCELL_36_352 ();
 FILLCELL_X32 FILLCELL_36_384 ();
 FILLCELL_X32 FILLCELL_36_416 ();
 FILLCELL_X32 FILLCELL_36_448 ();
 FILLCELL_X32 FILLCELL_36_480 ();
 FILLCELL_X32 FILLCELL_36_512 ();
 FILLCELL_X32 FILLCELL_36_544 ();
 FILLCELL_X32 FILLCELL_36_576 ();
 FILLCELL_X32 FILLCELL_36_608 ();
 FILLCELL_X32 FILLCELL_36_640 ();
 FILLCELL_X32 FILLCELL_36_672 ();
 FILLCELL_X32 FILLCELL_36_704 ();
 FILLCELL_X32 FILLCELL_36_736 ();
 FILLCELL_X32 FILLCELL_36_768 ();
 FILLCELL_X32 FILLCELL_36_800 ();
 FILLCELL_X32 FILLCELL_36_832 ();
 FILLCELL_X32 FILLCELL_36_864 ();
 FILLCELL_X32 FILLCELL_36_896 ();
 FILLCELL_X32 FILLCELL_36_928 ();
 FILLCELL_X32 FILLCELL_36_960 ();
 FILLCELL_X32 FILLCELL_36_992 ();
 FILLCELL_X32 FILLCELL_36_1024 ();
 FILLCELL_X32 FILLCELL_36_1056 ();
 FILLCELL_X32 FILLCELL_36_1088 ();
 FILLCELL_X32 FILLCELL_36_1120 ();
 FILLCELL_X32 FILLCELL_36_1152 ();
 FILLCELL_X32 FILLCELL_36_1184 ();
 FILLCELL_X32 FILLCELL_36_1216 ();
 FILLCELL_X32 FILLCELL_36_1248 ();
 FILLCELL_X32 FILLCELL_36_1280 ();
 FILLCELL_X32 FILLCELL_36_1312 ();
 FILLCELL_X32 FILLCELL_36_1344 ();
 FILLCELL_X32 FILLCELL_36_1376 ();
 FILLCELL_X32 FILLCELL_36_1408 ();
 FILLCELL_X32 FILLCELL_36_1440 ();
 FILLCELL_X32 FILLCELL_36_1472 ();
 FILLCELL_X32 FILLCELL_36_1504 ();
 FILLCELL_X32 FILLCELL_36_1536 ();
 FILLCELL_X32 FILLCELL_36_1568 ();
 FILLCELL_X32 FILLCELL_36_1600 ();
 FILLCELL_X32 FILLCELL_36_1632 ();
 FILLCELL_X32 FILLCELL_36_1664 ();
 FILLCELL_X32 FILLCELL_36_1696 ();
 FILLCELL_X32 FILLCELL_36_1728 ();
 FILLCELL_X32 FILLCELL_36_1760 ();
 FILLCELL_X32 FILLCELL_36_1792 ();
 FILLCELL_X32 FILLCELL_36_1824 ();
 FILLCELL_X32 FILLCELL_36_1856 ();
 FILLCELL_X8 FILLCELL_36_1888 ();
 FILLCELL_X1 FILLCELL_36_1896 ();
 FILLCELL_X32 FILLCELL_37_0 ();
 FILLCELL_X32 FILLCELL_37_32 ();
 FILLCELL_X32 FILLCELL_37_64 ();
 FILLCELL_X32 FILLCELL_37_96 ();
 FILLCELL_X32 FILLCELL_37_128 ();
 FILLCELL_X32 FILLCELL_37_160 ();
 FILLCELL_X32 FILLCELL_37_192 ();
 FILLCELL_X32 FILLCELL_37_224 ();
 FILLCELL_X32 FILLCELL_37_256 ();
 FILLCELL_X32 FILLCELL_37_288 ();
 FILLCELL_X32 FILLCELL_37_320 ();
 FILLCELL_X32 FILLCELL_37_352 ();
 FILLCELL_X32 FILLCELL_37_384 ();
 FILLCELL_X32 FILLCELL_37_416 ();
 FILLCELL_X32 FILLCELL_37_448 ();
 FILLCELL_X32 FILLCELL_37_480 ();
 FILLCELL_X32 FILLCELL_37_512 ();
 FILLCELL_X32 FILLCELL_37_544 ();
 FILLCELL_X32 FILLCELL_37_576 ();
 FILLCELL_X32 FILLCELL_37_608 ();
 FILLCELL_X32 FILLCELL_37_640 ();
 FILLCELL_X32 FILLCELL_37_672 ();
 FILLCELL_X32 FILLCELL_37_704 ();
 FILLCELL_X32 FILLCELL_37_736 ();
 FILLCELL_X32 FILLCELL_37_768 ();
 FILLCELL_X32 FILLCELL_37_800 ();
 FILLCELL_X32 FILLCELL_37_832 ();
 FILLCELL_X32 FILLCELL_37_864 ();
 FILLCELL_X32 FILLCELL_37_896 ();
 FILLCELL_X32 FILLCELL_37_928 ();
 FILLCELL_X32 FILLCELL_37_960 ();
 FILLCELL_X32 FILLCELL_37_992 ();
 FILLCELL_X32 FILLCELL_37_1024 ();
 FILLCELL_X32 FILLCELL_37_1056 ();
 FILLCELL_X32 FILLCELL_37_1088 ();
 FILLCELL_X32 FILLCELL_37_1120 ();
 FILLCELL_X32 FILLCELL_37_1152 ();
 FILLCELL_X32 FILLCELL_37_1184 ();
 FILLCELL_X32 FILLCELL_37_1216 ();
 FILLCELL_X32 FILLCELL_37_1248 ();
 FILLCELL_X32 FILLCELL_37_1280 ();
 FILLCELL_X32 FILLCELL_37_1312 ();
 FILLCELL_X32 FILLCELL_37_1344 ();
 FILLCELL_X32 FILLCELL_37_1376 ();
 FILLCELL_X32 FILLCELL_37_1408 ();
 FILLCELL_X32 FILLCELL_37_1440 ();
 FILLCELL_X32 FILLCELL_37_1472 ();
 FILLCELL_X32 FILLCELL_37_1504 ();
 FILLCELL_X32 FILLCELL_37_1536 ();
 FILLCELL_X32 FILLCELL_37_1568 ();
 FILLCELL_X32 FILLCELL_37_1600 ();
 FILLCELL_X32 FILLCELL_37_1632 ();
 FILLCELL_X32 FILLCELL_37_1664 ();
 FILLCELL_X32 FILLCELL_37_1696 ();
 FILLCELL_X32 FILLCELL_37_1728 ();
 FILLCELL_X32 FILLCELL_37_1760 ();
 FILLCELL_X32 FILLCELL_37_1792 ();
 FILLCELL_X32 FILLCELL_37_1824 ();
 FILLCELL_X32 FILLCELL_37_1856 ();
 FILLCELL_X8 FILLCELL_37_1888 ();
 FILLCELL_X1 FILLCELL_37_1896 ();
 FILLCELL_X32 FILLCELL_38_0 ();
 FILLCELL_X32 FILLCELL_38_32 ();
 FILLCELL_X32 FILLCELL_38_64 ();
 FILLCELL_X32 FILLCELL_38_96 ();
 FILLCELL_X32 FILLCELL_38_128 ();
 FILLCELL_X32 FILLCELL_38_160 ();
 FILLCELL_X32 FILLCELL_38_192 ();
 FILLCELL_X32 FILLCELL_38_224 ();
 FILLCELL_X32 FILLCELL_38_256 ();
 FILLCELL_X32 FILLCELL_38_288 ();
 FILLCELL_X32 FILLCELL_38_320 ();
 FILLCELL_X32 FILLCELL_38_352 ();
 FILLCELL_X32 FILLCELL_38_384 ();
 FILLCELL_X32 FILLCELL_38_416 ();
 FILLCELL_X32 FILLCELL_38_448 ();
 FILLCELL_X32 FILLCELL_38_480 ();
 FILLCELL_X32 FILLCELL_38_512 ();
 FILLCELL_X32 FILLCELL_38_544 ();
 FILLCELL_X32 FILLCELL_38_576 ();
 FILLCELL_X32 FILLCELL_38_608 ();
 FILLCELL_X32 FILLCELL_38_640 ();
 FILLCELL_X32 FILLCELL_38_672 ();
 FILLCELL_X32 FILLCELL_38_704 ();
 FILLCELL_X32 FILLCELL_38_736 ();
 FILLCELL_X32 FILLCELL_38_768 ();
 FILLCELL_X32 FILLCELL_38_800 ();
 FILLCELL_X32 FILLCELL_38_832 ();
 FILLCELL_X32 FILLCELL_38_864 ();
 FILLCELL_X32 FILLCELL_38_896 ();
 FILLCELL_X32 FILLCELL_38_928 ();
 FILLCELL_X32 FILLCELL_38_960 ();
 FILLCELL_X32 FILLCELL_38_992 ();
 FILLCELL_X32 FILLCELL_38_1024 ();
 FILLCELL_X32 FILLCELL_38_1056 ();
 FILLCELL_X32 FILLCELL_38_1088 ();
 FILLCELL_X32 FILLCELL_38_1120 ();
 FILLCELL_X32 FILLCELL_38_1152 ();
 FILLCELL_X32 FILLCELL_38_1184 ();
 FILLCELL_X32 FILLCELL_38_1216 ();
 FILLCELL_X32 FILLCELL_38_1248 ();
 FILLCELL_X32 FILLCELL_38_1280 ();
 FILLCELL_X32 FILLCELL_38_1312 ();
 FILLCELL_X32 FILLCELL_38_1344 ();
 FILLCELL_X32 FILLCELL_38_1376 ();
 FILLCELL_X32 FILLCELL_38_1408 ();
 FILLCELL_X32 FILLCELL_38_1440 ();
 FILLCELL_X32 FILLCELL_38_1472 ();
 FILLCELL_X32 FILLCELL_38_1504 ();
 FILLCELL_X32 FILLCELL_38_1536 ();
 FILLCELL_X32 FILLCELL_38_1568 ();
 FILLCELL_X32 FILLCELL_38_1600 ();
 FILLCELL_X32 FILLCELL_38_1632 ();
 FILLCELL_X32 FILLCELL_38_1664 ();
 FILLCELL_X32 FILLCELL_38_1696 ();
 FILLCELL_X32 FILLCELL_38_1728 ();
 FILLCELL_X32 FILLCELL_38_1760 ();
 FILLCELL_X32 FILLCELL_38_1792 ();
 FILLCELL_X32 FILLCELL_38_1824 ();
 FILLCELL_X32 FILLCELL_38_1856 ();
 FILLCELL_X8 FILLCELL_38_1888 ();
 FILLCELL_X1 FILLCELL_38_1896 ();
 FILLCELL_X32 FILLCELL_39_0 ();
 FILLCELL_X32 FILLCELL_39_32 ();
 FILLCELL_X32 FILLCELL_39_64 ();
 FILLCELL_X32 FILLCELL_39_96 ();
 FILLCELL_X32 FILLCELL_39_128 ();
 FILLCELL_X32 FILLCELL_39_160 ();
 FILLCELL_X32 FILLCELL_39_192 ();
 FILLCELL_X32 FILLCELL_39_224 ();
 FILLCELL_X32 FILLCELL_39_256 ();
 FILLCELL_X32 FILLCELL_39_288 ();
 FILLCELL_X32 FILLCELL_39_320 ();
 FILLCELL_X32 FILLCELL_39_352 ();
 FILLCELL_X32 FILLCELL_39_384 ();
 FILLCELL_X32 FILLCELL_39_416 ();
 FILLCELL_X32 FILLCELL_39_448 ();
 FILLCELL_X32 FILLCELL_39_480 ();
 FILLCELL_X32 FILLCELL_39_512 ();
 FILLCELL_X32 FILLCELL_39_544 ();
 FILLCELL_X32 FILLCELL_39_576 ();
 FILLCELL_X32 FILLCELL_39_608 ();
 FILLCELL_X32 FILLCELL_39_640 ();
 FILLCELL_X32 FILLCELL_39_672 ();
 FILLCELL_X32 FILLCELL_39_704 ();
 FILLCELL_X32 FILLCELL_39_736 ();
 FILLCELL_X32 FILLCELL_39_768 ();
 FILLCELL_X32 FILLCELL_39_800 ();
 FILLCELL_X32 FILLCELL_39_832 ();
 FILLCELL_X32 FILLCELL_39_864 ();
 FILLCELL_X32 FILLCELL_39_896 ();
 FILLCELL_X32 FILLCELL_39_928 ();
 FILLCELL_X32 FILLCELL_39_960 ();
 FILLCELL_X32 FILLCELL_39_992 ();
 FILLCELL_X32 FILLCELL_39_1024 ();
 FILLCELL_X32 FILLCELL_39_1056 ();
 FILLCELL_X32 FILLCELL_39_1088 ();
 FILLCELL_X32 FILLCELL_39_1120 ();
 FILLCELL_X32 FILLCELL_39_1152 ();
 FILLCELL_X32 FILLCELL_39_1184 ();
 FILLCELL_X32 FILLCELL_39_1216 ();
 FILLCELL_X32 FILLCELL_39_1248 ();
 FILLCELL_X32 FILLCELL_39_1280 ();
 FILLCELL_X32 FILLCELL_39_1312 ();
 FILLCELL_X32 FILLCELL_39_1344 ();
 FILLCELL_X32 FILLCELL_39_1376 ();
 FILLCELL_X32 FILLCELL_39_1408 ();
 FILLCELL_X32 FILLCELL_39_1440 ();
 FILLCELL_X32 FILLCELL_39_1472 ();
 FILLCELL_X32 FILLCELL_39_1504 ();
 FILLCELL_X32 FILLCELL_39_1536 ();
 FILLCELL_X32 FILLCELL_39_1568 ();
 FILLCELL_X32 FILLCELL_39_1600 ();
 FILLCELL_X32 FILLCELL_39_1632 ();
 FILLCELL_X32 FILLCELL_39_1664 ();
 FILLCELL_X32 FILLCELL_39_1696 ();
 FILLCELL_X32 FILLCELL_39_1728 ();
 FILLCELL_X32 FILLCELL_39_1760 ();
 FILLCELL_X32 FILLCELL_39_1792 ();
 FILLCELL_X32 FILLCELL_39_1824 ();
 FILLCELL_X32 FILLCELL_39_1856 ();
 FILLCELL_X8 FILLCELL_39_1888 ();
 FILLCELL_X1 FILLCELL_39_1896 ();
 FILLCELL_X32 FILLCELL_40_0 ();
 FILLCELL_X32 FILLCELL_40_32 ();
 FILLCELL_X32 FILLCELL_40_64 ();
 FILLCELL_X32 FILLCELL_40_96 ();
 FILLCELL_X32 FILLCELL_40_128 ();
 FILLCELL_X32 FILLCELL_40_160 ();
 FILLCELL_X32 FILLCELL_40_192 ();
 FILLCELL_X32 FILLCELL_40_224 ();
 FILLCELL_X32 FILLCELL_40_256 ();
 FILLCELL_X32 FILLCELL_40_288 ();
 FILLCELL_X32 FILLCELL_40_320 ();
 FILLCELL_X32 FILLCELL_40_352 ();
 FILLCELL_X32 FILLCELL_40_384 ();
 FILLCELL_X32 FILLCELL_40_416 ();
 FILLCELL_X32 FILLCELL_40_448 ();
 FILLCELL_X32 FILLCELL_40_480 ();
 FILLCELL_X32 FILLCELL_40_512 ();
 FILLCELL_X32 FILLCELL_40_544 ();
 FILLCELL_X32 FILLCELL_40_576 ();
 FILLCELL_X32 FILLCELL_40_608 ();
 FILLCELL_X32 FILLCELL_40_640 ();
 FILLCELL_X32 FILLCELL_40_672 ();
 FILLCELL_X32 FILLCELL_40_704 ();
 FILLCELL_X32 FILLCELL_40_736 ();
 FILLCELL_X32 FILLCELL_40_768 ();
 FILLCELL_X32 FILLCELL_40_800 ();
 FILLCELL_X32 FILLCELL_40_832 ();
 FILLCELL_X32 FILLCELL_40_864 ();
 FILLCELL_X32 FILLCELL_40_896 ();
 FILLCELL_X32 FILLCELL_40_928 ();
 FILLCELL_X32 FILLCELL_40_960 ();
 FILLCELL_X32 FILLCELL_40_992 ();
 FILLCELL_X32 FILLCELL_40_1024 ();
 FILLCELL_X32 FILLCELL_40_1056 ();
 FILLCELL_X32 FILLCELL_40_1088 ();
 FILLCELL_X32 FILLCELL_40_1120 ();
 FILLCELL_X32 FILLCELL_40_1152 ();
 FILLCELL_X32 FILLCELL_40_1184 ();
 FILLCELL_X32 FILLCELL_40_1216 ();
 FILLCELL_X32 FILLCELL_40_1248 ();
 FILLCELL_X32 FILLCELL_40_1280 ();
 FILLCELL_X32 FILLCELL_40_1312 ();
 FILLCELL_X32 FILLCELL_40_1344 ();
 FILLCELL_X32 FILLCELL_40_1376 ();
 FILLCELL_X32 FILLCELL_40_1408 ();
 FILLCELL_X32 FILLCELL_40_1440 ();
 FILLCELL_X32 FILLCELL_40_1472 ();
 FILLCELL_X32 FILLCELL_40_1504 ();
 FILLCELL_X32 FILLCELL_40_1536 ();
 FILLCELL_X32 FILLCELL_40_1568 ();
 FILLCELL_X32 FILLCELL_40_1600 ();
 FILLCELL_X32 FILLCELL_40_1632 ();
 FILLCELL_X32 FILLCELL_40_1664 ();
 FILLCELL_X32 FILLCELL_40_1696 ();
 FILLCELL_X32 FILLCELL_40_1728 ();
 FILLCELL_X32 FILLCELL_40_1760 ();
 FILLCELL_X32 FILLCELL_40_1792 ();
 FILLCELL_X32 FILLCELL_40_1824 ();
 FILLCELL_X32 FILLCELL_40_1856 ();
 FILLCELL_X8 FILLCELL_40_1888 ();
 FILLCELL_X1 FILLCELL_40_1896 ();
 FILLCELL_X32 FILLCELL_41_0 ();
 FILLCELL_X32 FILLCELL_41_32 ();
 FILLCELL_X32 FILLCELL_41_64 ();
 FILLCELL_X32 FILLCELL_41_96 ();
 FILLCELL_X32 FILLCELL_41_128 ();
 FILLCELL_X32 FILLCELL_41_160 ();
 FILLCELL_X32 FILLCELL_41_192 ();
 FILLCELL_X32 FILLCELL_41_224 ();
 FILLCELL_X32 FILLCELL_41_256 ();
 FILLCELL_X32 FILLCELL_41_288 ();
 FILLCELL_X32 FILLCELL_41_320 ();
 FILLCELL_X32 FILLCELL_41_352 ();
 FILLCELL_X32 FILLCELL_41_384 ();
 FILLCELL_X32 FILLCELL_41_416 ();
 FILLCELL_X32 FILLCELL_41_448 ();
 FILLCELL_X32 FILLCELL_41_480 ();
 FILLCELL_X32 FILLCELL_41_512 ();
 FILLCELL_X32 FILLCELL_41_544 ();
 FILLCELL_X32 FILLCELL_41_576 ();
 FILLCELL_X32 FILLCELL_41_608 ();
 FILLCELL_X32 FILLCELL_41_640 ();
 FILLCELL_X32 FILLCELL_41_672 ();
 FILLCELL_X32 FILLCELL_41_704 ();
 FILLCELL_X32 FILLCELL_41_736 ();
 FILLCELL_X32 FILLCELL_41_768 ();
 FILLCELL_X32 FILLCELL_41_800 ();
 FILLCELL_X32 FILLCELL_41_832 ();
 FILLCELL_X32 FILLCELL_41_864 ();
 FILLCELL_X32 FILLCELL_41_896 ();
 FILLCELL_X32 FILLCELL_41_928 ();
 FILLCELL_X32 FILLCELL_41_960 ();
 FILLCELL_X32 FILLCELL_41_992 ();
 FILLCELL_X32 FILLCELL_41_1024 ();
 FILLCELL_X32 FILLCELL_41_1056 ();
 FILLCELL_X32 FILLCELL_41_1088 ();
 FILLCELL_X32 FILLCELL_41_1120 ();
 FILLCELL_X32 FILLCELL_41_1152 ();
 FILLCELL_X32 FILLCELL_41_1184 ();
 FILLCELL_X32 FILLCELL_41_1216 ();
 FILLCELL_X32 FILLCELL_41_1248 ();
 FILLCELL_X32 FILLCELL_41_1280 ();
 FILLCELL_X32 FILLCELL_41_1312 ();
 FILLCELL_X32 FILLCELL_41_1344 ();
 FILLCELL_X32 FILLCELL_41_1376 ();
 FILLCELL_X32 FILLCELL_41_1408 ();
 FILLCELL_X32 FILLCELL_41_1440 ();
 FILLCELL_X32 FILLCELL_41_1472 ();
 FILLCELL_X32 FILLCELL_41_1504 ();
 FILLCELL_X32 FILLCELL_41_1536 ();
 FILLCELL_X32 FILLCELL_41_1568 ();
 FILLCELL_X32 FILLCELL_41_1600 ();
 FILLCELL_X32 FILLCELL_41_1632 ();
 FILLCELL_X32 FILLCELL_41_1664 ();
 FILLCELL_X32 FILLCELL_41_1696 ();
 FILLCELL_X32 FILLCELL_41_1728 ();
 FILLCELL_X32 FILLCELL_41_1760 ();
 FILLCELL_X32 FILLCELL_41_1792 ();
 FILLCELL_X32 FILLCELL_41_1824 ();
 FILLCELL_X32 FILLCELL_41_1856 ();
 FILLCELL_X8 FILLCELL_41_1888 ();
 FILLCELL_X1 FILLCELL_41_1896 ();
 FILLCELL_X32 FILLCELL_42_0 ();
 FILLCELL_X32 FILLCELL_42_32 ();
 FILLCELL_X32 FILLCELL_42_64 ();
 FILLCELL_X32 FILLCELL_42_96 ();
 FILLCELL_X32 FILLCELL_42_128 ();
 FILLCELL_X32 FILLCELL_42_160 ();
 FILLCELL_X32 FILLCELL_42_192 ();
 FILLCELL_X32 FILLCELL_42_224 ();
 FILLCELL_X32 FILLCELL_42_256 ();
 FILLCELL_X32 FILLCELL_42_288 ();
 FILLCELL_X32 FILLCELL_42_320 ();
 FILLCELL_X32 FILLCELL_42_352 ();
 FILLCELL_X32 FILLCELL_42_384 ();
 FILLCELL_X32 FILLCELL_42_416 ();
 FILLCELL_X32 FILLCELL_42_448 ();
 FILLCELL_X32 FILLCELL_42_480 ();
 FILLCELL_X32 FILLCELL_42_512 ();
 FILLCELL_X32 FILLCELL_42_544 ();
 FILLCELL_X32 FILLCELL_42_576 ();
 FILLCELL_X32 FILLCELL_42_608 ();
 FILLCELL_X32 FILLCELL_42_640 ();
 FILLCELL_X32 FILLCELL_42_672 ();
 FILLCELL_X32 FILLCELL_42_704 ();
 FILLCELL_X32 FILLCELL_42_736 ();
 FILLCELL_X32 FILLCELL_42_768 ();
 FILLCELL_X32 FILLCELL_42_800 ();
 FILLCELL_X32 FILLCELL_42_832 ();
 FILLCELL_X32 FILLCELL_42_864 ();
 FILLCELL_X32 FILLCELL_42_896 ();
 FILLCELL_X32 FILLCELL_42_928 ();
 FILLCELL_X32 FILLCELL_42_960 ();
 FILLCELL_X32 FILLCELL_42_992 ();
 FILLCELL_X32 FILLCELL_42_1024 ();
 FILLCELL_X32 FILLCELL_42_1056 ();
 FILLCELL_X32 FILLCELL_42_1088 ();
 FILLCELL_X32 FILLCELL_42_1120 ();
 FILLCELL_X32 FILLCELL_42_1152 ();
 FILLCELL_X32 FILLCELL_42_1184 ();
 FILLCELL_X32 FILLCELL_42_1216 ();
 FILLCELL_X32 FILLCELL_42_1248 ();
 FILLCELL_X32 FILLCELL_42_1280 ();
 FILLCELL_X32 FILLCELL_42_1312 ();
 FILLCELL_X32 FILLCELL_42_1344 ();
 FILLCELL_X32 FILLCELL_42_1376 ();
 FILLCELL_X32 FILLCELL_42_1408 ();
 FILLCELL_X32 FILLCELL_42_1440 ();
 FILLCELL_X32 FILLCELL_42_1472 ();
 FILLCELL_X32 FILLCELL_42_1504 ();
 FILLCELL_X32 FILLCELL_42_1536 ();
 FILLCELL_X32 FILLCELL_42_1568 ();
 FILLCELL_X32 FILLCELL_42_1600 ();
 FILLCELL_X32 FILLCELL_42_1632 ();
 FILLCELL_X32 FILLCELL_42_1664 ();
 FILLCELL_X32 FILLCELL_42_1696 ();
 FILLCELL_X32 FILLCELL_42_1728 ();
 FILLCELL_X32 FILLCELL_42_1760 ();
 FILLCELL_X32 FILLCELL_42_1792 ();
 FILLCELL_X32 FILLCELL_42_1824 ();
 FILLCELL_X32 FILLCELL_42_1856 ();
 FILLCELL_X8 FILLCELL_42_1888 ();
 FILLCELL_X1 FILLCELL_42_1896 ();
 FILLCELL_X32 FILLCELL_43_0 ();
 FILLCELL_X32 FILLCELL_43_32 ();
 FILLCELL_X32 FILLCELL_43_64 ();
 FILLCELL_X32 FILLCELL_43_96 ();
 FILLCELL_X32 FILLCELL_43_128 ();
 FILLCELL_X32 FILLCELL_43_160 ();
 FILLCELL_X32 FILLCELL_43_192 ();
 FILLCELL_X32 FILLCELL_43_224 ();
 FILLCELL_X32 FILLCELL_43_256 ();
 FILLCELL_X32 FILLCELL_43_288 ();
 FILLCELL_X32 FILLCELL_43_320 ();
 FILLCELL_X32 FILLCELL_43_352 ();
 FILLCELL_X32 FILLCELL_43_384 ();
 FILLCELL_X32 FILLCELL_43_416 ();
 FILLCELL_X32 FILLCELL_43_448 ();
 FILLCELL_X32 FILLCELL_43_480 ();
 FILLCELL_X32 FILLCELL_43_512 ();
 FILLCELL_X32 FILLCELL_43_544 ();
 FILLCELL_X32 FILLCELL_43_576 ();
 FILLCELL_X32 FILLCELL_43_608 ();
 FILLCELL_X32 FILLCELL_43_640 ();
 FILLCELL_X32 FILLCELL_43_672 ();
 FILLCELL_X32 FILLCELL_43_704 ();
 FILLCELL_X32 FILLCELL_43_736 ();
 FILLCELL_X32 FILLCELL_43_768 ();
 FILLCELL_X32 FILLCELL_43_800 ();
 FILLCELL_X32 FILLCELL_43_832 ();
 FILLCELL_X32 FILLCELL_43_864 ();
 FILLCELL_X32 FILLCELL_43_896 ();
 FILLCELL_X32 FILLCELL_43_928 ();
 FILLCELL_X32 FILLCELL_43_960 ();
 FILLCELL_X32 FILLCELL_43_992 ();
 FILLCELL_X32 FILLCELL_43_1024 ();
 FILLCELL_X32 FILLCELL_43_1056 ();
 FILLCELL_X32 FILLCELL_43_1088 ();
 FILLCELL_X32 FILLCELL_43_1120 ();
 FILLCELL_X32 FILLCELL_43_1152 ();
 FILLCELL_X32 FILLCELL_43_1184 ();
 FILLCELL_X32 FILLCELL_43_1216 ();
 FILLCELL_X32 FILLCELL_43_1248 ();
 FILLCELL_X32 FILLCELL_43_1280 ();
 FILLCELL_X32 FILLCELL_43_1312 ();
 FILLCELL_X32 FILLCELL_43_1344 ();
 FILLCELL_X32 FILLCELL_43_1376 ();
 FILLCELL_X32 FILLCELL_43_1408 ();
 FILLCELL_X32 FILLCELL_43_1440 ();
 FILLCELL_X32 FILLCELL_43_1472 ();
 FILLCELL_X32 FILLCELL_43_1504 ();
 FILLCELL_X32 FILLCELL_43_1536 ();
 FILLCELL_X32 FILLCELL_43_1568 ();
 FILLCELL_X32 FILLCELL_43_1600 ();
 FILLCELL_X32 FILLCELL_43_1632 ();
 FILLCELL_X32 FILLCELL_43_1664 ();
 FILLCELL_X32 FILLCELL_43_1696 ();
 FILLCELL_X32 FILLCELL_43_1728 ();
 FILLCELL_X32 FILLCELL_43_1760 ();
 FILLCELL_X32 FILLCELL_43_1792 ();
 FILLCELL_X32 FILLCELL_43_1824 ();
 FILLCELL_X32 FILLCELL_43_1856 ();
 FILLCELL_X8 FILLCELL_43_1888 ();
 FILLCELL_X1 FILLCELL_43_1896 ();
 FILLCELL_X32 FILLCELL_44_0 ();
 FILLCELL_X32 FILLCELL_44_32 ();
 FILLCELL_X32 FILLCELL_44_64 ();
 FILLCELL_X32 FILLCELL_44_96 ();
 FILLCELL_X32 FILLCELL_44_128 ();
 FILLCELL_X32 FILLCELL_44_160 ();
 FILLCELL_X32 FILLCELL_44_192 ();
 FILLCELL_X32 FILLCELL_44_224 ();
 FILLCELL_X32 FILLCELL_44_256 ();
 FILLCELL_X32 FILLCELL_44_288 ();
 FILLCELL_X32 FILLCELL_44_320 ();
 FILLCELL_X32 FILLCELL_44_352 ();
 FILLCELL_X32 FILLCELL_44_384 ();
 FILLCELL_X32 FILLCELL_44_416 ();
 FILLCELL_X32 FILLCELL_44_448 ();
 FILLCELL_X32 FILLCELL_44_480 ();
 FILLCELL_X32 FILLCELL_44_512 ();
 FILLCELL_X32 FILLCELL_44_544 ();
 FILLCELL_X32 FILLCELL_44_576 ();
 FILLCELL_X32 FILLCELL_44_608 ();
 FILLCELL_X32 FILLCELL_44_640 ();
 FILLCELL_X32 FILLCELL_44_672 ();
 FILLCELL_X32 FILLCELL_44_704 ();
 FILLCELL_X32 FILLCELL_44_736 ();
 FILLCELL_X32 FILLCELL_44_768 ();
 FILLCELL_X32 FILLCELL_44_800 ();
 FILLCELL_X32 FILLCELL_44_832 ();
 FILLCELL_X32 FILLCELL_44_864 ();
 FILLCELL_X32 FILLCELL_44_896 ();
 FILLCELL_X32 FILLCELL_44_928 ();
 FILLCELL_X32 FILLCELL_44_960 ();
 FILLCELL_X32 FILLCELL_44_992 ();
 FILLCELL_X32 FILLCELL_44_1024 ();
 FILLCELL_X32 FILLCELL_44_1056 ();
 FILLCELL_X32 FILLCELL_44_1088 ();
 FILLCELL_X32 FILLCELL_44_1120 ();
 FILLCELL_X32 FILLCELL_44_1152 ();
 FILLCELL_X32 FILLCELL_44_1184 ();
 FILLCELL_X32 FILLCELL_44_1216 ();
 FILLCELL_X32 FILLCELL_44_1248 ();
 FILLCELL_X32 FILLCELL_44_1280 ();
 FILLCELL_X32 FILLCELL_44_1312 ();
 FILLCELL_X32 FILLCELL_44_1344 ();
 FILLCELL_X32 FILLCELL_44_1376 ();
 FILLCELL_X32 FILLCELL_44_1408 ();
 FILLCELL_X32 FILLCELL_44_1440 ();
 FILLCELL_X32 FILLCELL_44_1472 ();
 FILLCELL_X32 FILLCELL_44_1504 ();
 FILLCELL_X32 FILLCELL_44_1536 ();
 FILLCELL_X32 FILLCELL_44_1568 ();
 FILLCELL_X32 FILLCELL_44_1600 ();
 FILLCELL_X32 FILLCELL_44_1632 ();
 FILLCELL_X32 FILLCELL_44_1664 ();
 FILLCELL_X32 FILLCELL_44_1696 ();
 FILLCELL_X32 FILLCELL_44_1728 ();
 FILLCELL_X32 FILLCELL_44_1760 ();
 FILLCELL_X32 FILLCELL_44_1792 ();
 FILLCELL_X32 FILLCELL_44_1824 ();
 FILLCELL_X32 FILLCELL_44_1856 ();
 FILLCELL_X8 FILLCELL_44_1888 ();
 FILLCELL_X1 FILLCELL_44_1896 ();
 FILLCELL_X32 FILLCELL_45_0 ();
 FILLCELL_X32 FILLCELL_45_32 ();
 FILLCELL_X32 FILLCELL_45_64 ();
 FILLCELL_X32 FILLCELL_45_96 ();
 FILLCELL_X32 FILLCELL_45_128 ();
 FILLCELL_X32 FILLCELL_45_160 ();
 FILLCELL_X32 FILLCELL_45_192 ();
 FILLCELL_X32 FILLCELL_45_224 ();
 FILLCELL_X32 FILLCELL_45_256 ();
 FILLCELL_X32 FILLCELL_45_288 ();
 FILLCELL_X32 FILLCELL_45_320 ();
 FILLCELL_X32 FILLCELL_45_352 ();
 FILLCELL_X32 FILLCELL_45_384 ();
 FILLCELL_X32 FILLCELL_45_416 ();
 FILLCELL_X32 FILLCELL_45_448 ();
 FILLCELL_X32 FILLCELL_45_480 ();
 FILLCELL_X32 FILLCELL_45_512 ();
 FILLCELL_X32 FILLCELL_45_544 ();
 FILLCELL_X32 FILLCELL_45_576 ();
 FILLCELL_X32 FILLCELL_45_608 ();
 FILLCELL_X32 FILLCELL_45_640 ();
 FILLCELL_X32 FILLCELL_45_672 ();
 FILLCELL_X32 FILLCELL_45_704 ();
 FILLCELL_X32 FILLCELL_45_736 ();
 FILLCELL_X32 FILLCELL_45_768 ();
 FILLCELL_X32 FILLCELL_45_800 ();
 FILLCELL_X32 FILLCELL_45_832 ();
 FILLCELL_X32 FILLCELL_45_864 ();
 FILLCELL_X32 FILLCELL_45_896 ();
 FILLCELL_X32 FILLCELL_45_928 ();
 FILLCELL_X32 FILLCELL_45_960 ();
 FILLCELL_X32 FILLCELL_45_992 ();
 FILLCELL_X32 FILLCELL_45_1024 ();
 FILLCELL_X32 FILLCELL_45_1056 ();
 FILLCELL_X32 FILLCELL_45_1088 ();
 FILLCELL_X32 FILLCELL_45_1120 ();
 FILLCELL_X32 FILLCELL_45_1152 ();
 FILLCELL_X32 FILLCELL_45_1184 ();
 FILLCELL_X32 FILLCELL_45_1216 ();
 FILLCELL_X32 FILLCELL_45_1248 ();
 FILLCELL_X32 FILLCELL_45_1280 ();
 FILLCELL_X32 FILLCELL_45_1312 ();
 FILLCELL_X32 FILLCELL_45_1344 ();
 FILLCELL_X32 FILLCELL_45_1376 ();
 FILLCELL_X32 FILLCELL_45_1408 ();
 FILLCELL_X32 FILLCELL_45_1440 ();
 FILLCELL_X32 FILLCELL_45_1472 ();
 FILLCELL_X32 FILLCELL_45_1504 ();
 FILLCELL_X32 FILLCELL_45_1536 ();
 FILLCELL_X32 FILLCELL_45_1568 ();
 FILLCELL_X32 FILLCELL_45_1600 ();
 FILLCELL_X32 FILLCELL_45_1632 ();
 FILLCELL_X32 FILLCELL_45_1664 ();
 FILLCELL_X32 FILLCELL_45_1696 ();
 FILLCELL_X32 FILLCELL_45_1728 ();
 FILLCELL_X32 FILLCELL_45_1760 ();
 FILLCELL_X32 FILLCELL_45_1792 ();
 FILLCELL_X32 FILLCELL_45_1824 ();
 FILLCELL_X32 FILLCELL_45_1856 ();
 FILLCELL_X8 FILLCELL_45_1888 ();
 FILLCELL_X1 FILLCELL_45_1896 ();
 FILLCELL_X32 FILLCELL_46_0 ();
 FILLCELL_X32 FILLCELL_46_32 ();
 FILLCELL_X32 FILLCELL_46_64 ();
 FILLCELL_X32 FILLCELL_46_96 ();
 FILLCELL_X32 FILLCELL_46_128 ();
 FILLCELL_X32 FILLCELL_46_160 ();
 FILLCELL_X32 FILLCELL_46_192 ();
 FILLCELL_X32 FILLCELL_46_224 ();
 FILLCELL_X32 FILLCELL_46_256 ();
 FILLCELL_X32 FILLCELL_46_288 ();
 FILLCELL_X32 FILLCELL_46_320 ();
 FILLCELL_X32 FILLCELL_46_352 ();
 FILLCELL_X32 FILLCELL_46_384 ();
 FILLCELL_X32 FILLCELL_46_416 ();
 FILLCELL_X32 FILLCELL_46_448 ();
 FILLCELL_X32 FILLCELL_46_480 ();
 FILLCELL_X32 FILLCELL_46_512 ();
 FILLCELL_X32 FILLCELL_46_544 ();
 FILLCELL_X32 FILLCELL_46_576 ();
 FILLCELL_X32 FILLCELL_46_608 ();
 FILLCELL_X32 FILLCELL_46_640 ();
 FILLCELL_X32 FILLCELL_46_672 ();
 FILLCELL_X32 FILLCELL_46_704 ();
 FILLCELL_X32 FILLCELL_46_736 ();
 FILLCELL_X32 FILLCELL_46_768 ();
 FILLCELL_X32 FILLCELL_46_800 ();
 FILLCELL_X32 FILLCELL_46_832 ();
 FILLCELL_X32 FILLCELL_46_864 ();
 FILLCELL_X32 FILLCELL_46_896 ();
 FILLCELL_X32 FILLCELL_46_928 ();
 FILLCELL_X32 FILLCELL_46_960 ();
 FILLCELL_X32 FILLCELL_46_992 ();
 FILLCELL_X32 FILLCELL_46_1024 ();
 FILLCELL_X32 FILLCELL_46_1056 ();
 FILLCELL_X32 FILLCELL_46_1088 ();
 FILLCELL_X32 FILLCELL_46_1120 ();
 FILLCELL_X32 FILLCELL_46_1152 ();
 FILLCELL_X32 FILLCELL_46_1184 ();
 FILLCELL_X32 FILLCELL_46_1216 ();
 FILLCELL_X32 FILLCELL_46_1248 ();
 FILLCELL_X32 FILLCELL_46_1280 ();
 FILLCELL_X32 FILLCELL_46_1312 ();
 FILLCELL_X32 FILLCELL_46_1344 ();
 FILLCELL_X32 FILLCELL_46_1376 ();
 FILLCELL_X32 FILLCELL_46_1408 ();
 FILLCELL_X32 FILLCELL_46_1440 ();
 FILLCELL_X32 FILLCELL_46_1472 ();
 FILLCELL_X32 FILLCELL_46_1504 ();
 FILLCELL_X32 FILLCELL_46_1536 ();
 FILLCELL_X32 FILLCELL_46_1568 ();
 FILLCELL_X32 FILLCELL_46_1600 ();
 FILLCELL_X32 FILLCELL_46_1632 ();
 FILLCELL_X32 FILLCELL_46_1664 ();
 FILLCELL_X32 FILLCELL_46_1696 ();
 FILLCELL_X32 FILLCELL_46_1728 ();
 FILLCELL_X32 FILLCELL_46_1760 ();
 FILLCELL_X32 FILLCELL_46_1792 ();
 FILLCELL_X32 FILLCELL_46_1824 ();
 FILLCELL_X32 FILLCELL_46_1856 ();
 FILLCELL_X8 FILLCELL_46_1888 ();
 FILLCELL_X1 FILLCELL_46_1896 ();
 FILLCELL_X32 FILLCELL_47_0 ();
 FILLCELL_X32 FILLCELL_47_32 ();
 FILLCELL_X32 FILLCELL_47_64 ();
 FILLCELL_X32 FILLCELL_47_96 ();
 FILLCELL_X32 FILLCELL_47_128 ();
 FILLCELL_X32 FILLCELL_47_160 ();
 FILLCELL_X32 FILLCELL_47_192 ();
 FILLCELL_X32 FILLCELL_47_224 ();
 FILLCELL_X32 FILLCELL_47_256 ();
 FILLCELL_X32 FILLCELL_47_288 ();
 FILLCELL_X32 FILLCELL_47_320 ();
 FILLCELL_X32 FILLCELL_47_352 ();
 FILLCELL_X32 FILLCELL_47_384 ();
 FILLCELL_X32 FILLCELL_47_416 ();
 FILLCELL_X32 FILLCELL_47_448 ();
 FILLCELL_X32 FILLCELL_47_480 ();
 FILLCELL_X32 FILLCELL_47_512 ();
 FILLCELL_X32 FILLCELL_47_544 ();
 FILLCELL_X32 FILLCELL_47_576 ();
 FILLCELL_X32 FILLCELL_47_608 ();
 FILLCELL_X32 FILLCELL_47_640 ();
 FILLCELL_X32 FILLCELL_47_672 ();
 FILLCELL_X32 FILLCELL_47_704 ();
 FILLCELL_X32 FILLCELL_47_736 ();
 FILLCELL_X32 FILLCELL_47_768 ();
 FILLCELL_X32 FILLCELL_47_800 ();
 FILLCELL_X32 FILLCELL_47_832 ();
 FILLCELL_X32 FILLCELL_47_864 ();
 FILLCELL_X32 FILLCELL_47_896 ();
 FILLCELL_X32 FILLCELL_47_928 ();
 FILLCELL_X32 FILLCELL_47_960 ();
 FILLCELL_X32 FILLCELL_47_992 ();
 FILLCELL_X32 FILLCELL_47_1024 ();
 FILLCELL_X32 FILLCELL_47_1056 ();
 FILLCELL_X32 FILLCELL_47_1088 ();
 FILLCELL_X32 FILLCELL_47_1120 ();
 FILLCELL_X32 FILLCELL_47_1152 ();
 FILLCELL_X32 FILLCELL_47_1184 ();
 FILLCELL_X32 FILLCELL_47_1216 ();
 FILLCELL_X32 FILLCELL_47_1248 ();
 FILLCELL_X32 FILLCELL_47_1280 ();
 FILLCELL_X32 FILLCELL_47_1312 ();
 FILLCELL_X32 FILLCELL_47_1344 ();
 FILLCELL_X32 FILLCELL_47_1376 ();
 FILLCELL_X32 FILLCELL_47_1408 ();
 FILLCELL_X32 FILLCELL_47_1440 ();
 FILLCELL_X32 FILLCELL_47_1472 ();
 FILLCELL_X32 FILLCELL_47_1504 ();
 FILLCELL_X32 FILLCELL_47_1536 ();
 FILLCELL_X32 FILLCELL_47_1568 ();
 FILLCELL_X32 FILLCELL_47_1600 ();
 FILLCELL_X32 FILLCELL_47_1632 ();
 FILLCELL_X32 FILLCELL_47_1664 ();
 FILLCELL_X32 FILLCELL_47_1696 ();
 FILLCELL_X32 FILLCELL_47_1728 ();
 FILLCELL_X32 FILLCELL_47_1760 ();
 FILLCELL_X32 FILLCELL_47_1792 ();
 FILLCELL_X32 FILLCELL_47_1824 ();
 FILLCELL_X32 FILLCELL_47_1856 ();
 FILLCELL_X8 FILLCELL_47_1888 ();
 FILLCELL_X1 FILLCELL_47_1896 ();
 FILLCELL_X32 FILLCELL_48_0 ();
 FILLCELL_X32 FILLCELL_48_32 ();
 FILLCELL_X32 FILLCELL_48_64 ();
 FILLCELL_X32 FILLCELL_48_96 ();
 FILLCELL_X32 FILLCELL_48_128 ();
 FILLCELL_X32 FILLCELL_48_160 ();
 FILLCELL_X32 FILLCELL_48_192 ();
 FILLCELL_X32 FILLCELL_48_224 ();
 FILLCELL_X32 FILLCELL_48_256 ();
 FILLCELL_X32 FILLCELL_48_288 ();
 FILLCELL_X32 FILLCELL_48_320 ();
 FILLCELL_X32 FILLCELL_48_352 ();
 FILLCELL_X32 FILLCELL_48_384 ();
 FILLCELL_X32 FILLCELL_48_416 ();
 FILLCELL_X32 FILLCELL_48_448 ();
 FILLCELL_X32 FILLCELL_48_480 ();
 FILLCELL_X32 FILLCELL_48_512 ();
 FILLCELL_X32 FILLCELL_48_544 ();
 FILLCELL_X32 FILLCELL_48_576 ();
 FILLCELL_X32 FILLCELL_48_608 ();
 FILLCELL_X32 FILLCELL_48_640 ();
 FILLCELL_X32 FILLCELL_48_672 ();
 FILLCELL_X32 FILLCELL_48_704 ();
 FILLCELL_X32 FILLCELL_48_736 ();
 FILLCELL_X32 FILLCELL_48_768 ();
 FILLCELL_X32 FILLCELL_48_800 ();
 FILLCELL_X32 FILLCELL_48_832 ();
 FILLCELL_X32 FILLCELL_48_864 ();
 FILLCELL_X32 FILLCELL_48_896 ();
 FILLCELL_X32 FILLCELL_48_928 ();
 FILLCELL_X32 FILLCELL_48_960 ();
 FILLCELL_X32 FILLCELL_48_992 ();
 FILLCELL_X32 FILLCELL_48_1024 ();
 FILLCELL_X32 FILLCELL_48_1056 ();
 FILLCELL_X32 FILLCELL_48_1088 ();
 FILLCELL_X32 FILLCELL_48_1120 ();
 FILLCELL_X32 FILLCELL_48_1152 ();
 FILLCELL_X32 FILLCELL_48_1184 ();
 FILLCELL_X32 FILLCELL_48_1216 ();
 FILLCELL_X32 FILLCELL_48_1248 ();
 FILLCELL_X32 FILLCELL_48_1280 ();
 FILLCELL_X32 FILLCELL_48_1312 ();
 FILLCELL_X32 FILLCELL_48_1344 ();
 FILLCELL_X32 FILLCELL_48_1376 ();
 FILLCELL_X32 FILLCELL_48_1408 ();
 FILLCELL_X32 FILLCELL_48_1440 ();
 FILLCELL_X32 FILLCELL_48_1472 ();
 FILLCELL_X32 FILLCELL_48_1504 ();
 FILLCELL_X32 FILLCELL_48_1536 ();
 FILLCELL_X32 FILLCELL_48_1568 ();
 FILLCELL_X32 FILLCELL_48_1600 ();
 FILLCELL_X32 FILLCELL_48_1632 ();
 FILLCELL_X32 FILLCELL_48_1664 ();
 FILLCELL_X32 FILLCELL_48_1696 ();
 FILLCELL_X32 FILLCELL_48_1728 ();
 FILLCELL_X32 FILLCELL_48_1760 ();
 FILLCELL_X32 FILLCELL_48_1792 ();
 FILLCELL_X32 FILLCELL_48_1824 ();
 FILLCELL_X32 FILLCELL_48_1856 ();
 FILLCELL_X8 FILLCELL_48_1888 ();
 FILLCELL_X1 FILLCELL_48_1896 ();
 FILLCELL_X32 FILLCELL_49_0 ();
 FILLCELL_X32 FILLCELL_49_32 ();
 FILLCELL_X32 FILLCELL_49_64 ();
 FILLCELL_X32 FILLCELL_49_96 ();
 FILLCELL_X32 FILLCELL_49_128 ();
 FILLCELL_X32 FILLCELL_49_160 ();
 FILLCELL_X32 FILLCELL_49_192 ();
 FILLCELL_X32 FILLCELL_49_224 ();
 FILLCELL_X32 FILLCELL_49_256 ();
 FILLCELL_X32 FILLCELL_49_288 ();
 FILLCELL_X32 FILLCELL_49_320 ();
 FILLCELL_X32 FILLCELL_49_352 ();
 FILLCELL_X32 FILLCELL_49_384 ();
 FILLCELL_X32 FILLCELL_49_416 ();
 FILLCELL_X32 FILLCELL_49_448 ();
 FILLCELL_X32 FILLCELL_49_480 ();
 FILLCELL_X32 FILLCELL_49_512 ();
 FILLCELL_X32 FILLCELL_49_544 ();
 FILLCELL_X32 FILLCELL_49_576 ();
 FILLCELL_X32 FILLCELL_49_608 ();
 FILLCELL_X32 FILLCELL_49_640 ();
 FILLCELL_X32 FILLCELL_49_672 ();
 FILLCELL_X32 FILLCELL_49_704 ();
 FILLCELL_X32 FILLCELL_49_736 ();
 FILLCELL_X32 FILLCELL_49_768 ();
 FILLCELL_X32 FILLCELL_49_800 ();
 FILLCELL_X32 FILLCELL_49_832 ();
 FILLCELL_X32 FILLCELL_49_864 ();
 FILLCELL_X32 FILLCELL_49_896 ();
 FILLCELL_X32 FILLCELL_49_928 ();
 FILLCELL_X32 FILLCELL_49_960 ();
 FILLCELL_X32 FILLCELL_49_992 ();
 FILLCELL_X32 FILLCELL_49_1024 ();
 FILLCELL_X32 FILLCELL_49_1056 ();
 FILLCELL_X32 FILLCELL_49_1088 ();
 FILLCELL_X32 FILLCELL_49_1120 ();
 FILLCELL_X32 FILLCELL_49_1152 ();
 FILLCELL_X32 FILLCELL_49_1184 ();
 FILLCELL_X32 FILLCELL_49_1216 ();
 FILLCELL_X32 FILLCELL_49_1248 ();
 FILLCELL_X32 FILLCELL_49_1280 ();
 FILLCELL_X32 FILLCELL_49_1312 ();
 FILLCELL_X32 FILLCELL_49_1344 ();
 FILLCELL_X32 FILLCELL_49_1376 ();
 FILLCELL_X32 FILLCELL_49_1408 ();
 FILLCELL_X32 FILLCELL_49_1440 ();
 FILLCELL_X32 FILLCELL_49_1472 ();
 FILLCELL_X32 FILLCELL_49_1504 ();
 FILLCELL_X32 FILLCELL_49_1536 ();
 FILLCELL_X32 FILLCELL_49_1568 ();
 FILLCELL_X32 FILLCELL_49_1600 ();
 FILLCELL_X32 FILLCELL_49_1632 ();
 FILLCELL_X32 FILLCELL_49_1664 ();
 FILLCELL_X32 FILLCELL_49_1696 ();
 FILLCELL_X32 FILLCELL_49_1728 ();
 FILLCELL_X32 FILLCELL_49_1760 ();
 FILLCELL_X32 FILLCELL_49_1792 ();
 FILLCELL_X32 FILLCELL_49_1824 ();
 FILLCELL_X32 FILLCELL_49_1856 ();
 FILLCELL_X8 FILLCELL_49_1888 ();
 FILLCELL_X1 FILLCELL_49_1896 ();
 FILLCELL_X32 FILLCELL_50_0 ();
 FILLCELL_X32 FILLCELL_50_32 ();
 FILLCELL_X32 FILLCELL_50_64 ();
 FILLCELL_X32 FILLCELL_50_96 ();
 FILLCELL_X32 FILLCELL_50_128 ();
 FILLCELL_X32 FILLCELL_50_160 ();
 FILLCELL_X32 FILLCELL_50_192 ();
 FILLCELL_X32 FILLCELL_50_224 ();
 FILLCELL_X32 FILLCELL_50_256 ();
 FILLCELL_X32 FILLCELL_50_288 ();
 FILLCELL_X32 FILLCELL_50_320 ();
 FILLCELL_X32 FILLCELL_50_352 ();
 FILLCELL_X32 FILLCELL_50_384 ();
 FILLCELL_X32 FILLCELL_50_416 ();
 FILLCELL_X32 FILLCELL_50_448 ();
 FILLCELL_X32 FILLCELL_50_480 ();
 FILLCELL_X32 FILLCELL_50_512 ();
 FILLCELL_X32 FILLCELL_50_544 ();
 FILLCELL_X32 FILLCELL_50_576 ();
 FILLCELL_X32 FILLCELL_50_608 ();
 FILLCELL_X32 FILLCELL_50_640 ();
 FILLCELL_X32 FILLCELL_50_672 ();
 FILLCELL_X32 FILLCELL_50_704 ();
 FILLCELL_X32 FILLCELL_50_736 ();
 FILLCELL_X32 FILLCELL_50_768 ();
 FILLCELL_X32 FILLCELL_50_800 ();
 FILLCELL_X32 FILLCELL_50_832 ();
 FILLCELL_X32 FILLCELL_50_864 ();
 FILLCELL_X32 FILLCELL_50_896 ();
 FILLCELL_X32 FILLCELL_50_928 ();
 FILLCELL_X32 FILLCELL_50_960 ();
 FILLCELL_X32 FILLCELL_50_992 ();
 FILLCELL_X32 FILLCELL_50_1024 ();
 FILLCELL_X32 FILLCELL_50_1056 ();
 FILLCELL_X32 FILLCELL_50_1088 ();
 FILLCELL_X32 FILLCELL_50_1120 ();
 FILLCELL_X32 FILLCELL_50_1152 ();
 FILLCELL_X32 FILLCELL_50_1184 ();
 FILLCELL_X32 FILLCELL_50_1216 ();
 FILLCELL_X32 FILLCELL_50_1248 ();
 FILLCELL_X32 FILLCELL_50_1280 ();
 FILLCELL_X32 FILLCELL_50_1312 ();
 FILLCELL_X32 FILLCELL_50_1344 ();
 FILLCELL_X32 FILLCELL_50_1376 ();
 FILLCELL_X32 FILLCELL_50_1408 ();
 FILLCELL_X32 FILLCELL_50_1440 ();
 FILLCELL_X32 FILLCELL_50_1472 ();
 FILLCELL_X32 FILLCELL_50_1504 ();
 FILLCELL_X32 FILLCELL_50_1536 ();
 FILLCELL_X32 FILLCELL_50_1568 ();
 FILLCELL_X32 FILLCELL_50_1600 ();
 FILLCELL_X32 FILLCELL_50_1632 ();
 FILLCELL_X32 FILLCELL_50_1664 ();
 FILLCELL_X32 FILLCELL_50_1696 ();
 FILLCELL_X32 FILLCELL_50_1728 ();
 FILLCELL_X32 FILLCELL_50_1760 ();
 FILLCELL_X32 FILLCELL_50_1792 ();
 FILLCELL_X32 FILLCELL_50_1824 ();
 FILLCELL_X32 FILLCELL_50_1856 ();
 FILLCELL_X8 FILLCELL_50_1888 ();
 FILLCELL_X1 FILLCELL_50_1896 ();
 FILLCELL_X32 FILLCELL_51_0 ();
 FILLCELL_X32 FILLCELL_51_32 ();
 FILLCELL_X32 FILLCELL_51_64 ();
 FILLCELL_X32 FILLCELL_51_96 ();
 FILLCELL_X32 FILLCELL_51_128 ();
 FILLCELL_X32 FILLCELL_51_160 ();
 FILLCELL_X32 FILLCELL_51_192 ();
 FILLCELL_X32 FILLCELL_51_224 ();
 FILLCELL_X32 FILLCELL_51_256 ();
 FILLCELL_X32 FILLCELL_51_288 ();
 FILLCELL_X32 FILLCELL_51_320 ();
 FILLCELL_X32 FILLCELL_51_352 ();
 FILLCELL_X32 FILLCELL_51_384 ();
 FILLCELL_X32 FILLCELL_51_416 ();
 FILLCELL_X32 FILLCELL_51_448 ();
 FILLCELL_X32 FILLCELL_51_480 ();
 FILLCELL_X32 FILLCELL_51_512 ();
 FILLCELL_X32 FILLCELL_51_544 ();
 FILLCELL_X32 FILLCELL_51_576 ();
 FILLCELL_X32 FILLCELL_51_608 ();
 FILLCELL_X32 FILLCELL_51_640 ();
 FILLCELL_X32 FILLCELL_51_672 ();
 FILLCELL_X32 FILLCELL_51_704 ();
 FILLCELL_X32 FILLCELL_51_736 ();
 FILLCELL_X32 FILLCELL_51_768 ();
 FILLCELL_X32 FILLCELL_51_800 ();
 FILLCELL_X32 FILLCELL_51_832 ();
 FILLCELL_X32 FILLCELL_51_864 ();
 FILLCELL_X32 FILLCELL_51_896 ();
 FILLCELL_X32 FILLCELL_51_928 ();
 FILLCELL_X32 FILLCELL_51_960 ();
 FILLCELL_X32 FILLCELL_51_992 ();
 FILLCELL_X32 FILLCELL_51_1024 ();
 FILLCELL_X32 FILLCELL_51_1056 ();
 FILLCELL_X32 FILLCELL_51_1088 ();
 FILLCELL_X32 FILLCELL_51_1120 ();
 FILLCELL_X32 FILLCELL_51_1152 ();
 FILLCELL_X32 FILLCELL_51_1184 ();
 FILLCELL_X32 FILLCELL_51_1216 ();
 FILLCELL_X32 FILLCELL_51_1248 ();
 FILLCELL_X32 FILLCELL_51_1280 ();
 FILLCELL_X32 FILLCELL_51_1312 ();
 FILLCELL_X32 FILLCELL_51_1344 ();
 FILLCELL_X32 FILLCELL_51_1376 ();
 FILLCELL_X32 FILLCELL_51_1408 ();
 FILLCELL_X32 FILLCELL_51_1440 ();
 FILLCELL_X32 FILLCELL_51_1472 ();
 FILLCELL_X32 FILLCELL_51_1504 ();
 FILLCELL_X32 FILLCELL_51_1536 ();
 FILLCELL_X32 FILLCELL_51_1568 ();
 FILLCELL_X32 FILLCELL_51_1600 ();
 FILLCELL_X32 FILLCELL_51_1632 ();
 FILLCELL_X32 FILLCELL_51_1664 ();
 FILLCELL_X32 FILLCELL_51_1696 ();
 FILLCELL_X32 FILLCELL_51_1728 ();
 FILLCELL_X32 FILLCELL_51_1760 ();
 FILLCELL_X32 FILLCELL_51_1792 ();
 FILLCELL_X32 FILLCELL_51_1824 ();
 FILLCELL_X32 FILLCELL_51_1856 ();
 FILLCELL_X8 FILLCELL_51_1888 ();
 FILLCELL_X1 FILLCELL_51_1896 ();
 FILLCELL_X32 FILLCELL_52_0 ();
 FILLCELL_X32 FILLCELL_52_32 ();
 FILLCELL_X32 FILLCELL_52_64 ();
 FILLCELL_X32 FILLCELL_52_96 ();
 FILLCELL_X32 FILLCELL_52_128 ();
 FILLCELL_X32 FILLCELL_52_160 ();
 FILLCELL_X32 FILLCELL_52_192 ();
 FILLCELL_X32 FILLCELL_52_224 ();
 FILLCELL_X32 FILLCELL_52_256 ();
 FILLCELL_X32 FILLCELL_52_288 ();
 FILLCELL_X32 FILLCELL_52_320 ();
 FILLCELL_X32 FILLCELL_52_352 ();
 FILLCELL_X32 FILLCELL_52_384 ();
 FILLCELL_X32 FILLCELL_52_416 ();
 FILLCELL_X16 FILLCELL_52_448 ();
 FILLCELL_X8 FILLCELL_52_464 ();
 FILLCELL_X4 FILLCELL_52_472 ();
 FILLCELL_X2 FILLCELL_52_476 ();
 FILLCELL_X32 FILLCELL_52_495 ();
 FILLCELL_X32 FILLCELL_52_527 ();
 FILLCELL_X32 FILLCELL_52_559 ();
 FILLCELL_X32 FILLCELL_52_591 ();
 FILLCELL_X32 FILLCELL_52_623 ();
 FILLCELL_X32 FILLCELL_52_655 ();
 FILLCELL_X32 FILLCELL_52_687 ();
 FILLCELL_X32 FILLCELL_52_719 ();
 FILLCELL_X32 FILLCELL_52_751 ();
 FILLCELL_X32 FILLCELL_52_783 ();
 FILLCELL_X32 FILLCELL_52_815 ();
 FILLCELL_X32 FILLCELL_52_847 ();
 FILLCELL_X32 FILLCELL_52_879 ();
 FILLCELL_X32 FILLCELL_52_911 ();
 FILLCELL_X32 FILLCELL_52_943 ();
 FILLCELL_X32 FILLCELL_52_975 ();
 FILLCELL_X32 FILLCELL_52_1007 ();
 FILLCELL_X32 FILLCELL_52_1039 ();
 FILLCELL_X32 FILLCELL_52_1071 ();
 FILLCELL_X32 FILLCELL_52_1103 ();
 FILLCELL_X32 FILLCELL_52_1135 ();
 FILLCELL_X32 FILLCELL_52_1167 ();
 FILLCELL_X32 FILLCELL_52_1199 ();
 FILLCELL_X32 FILLCELL_52_1231 ();
 FILLCELL_X32 FILLCELL_52_1263 ();
 FILLCELL_X32 FILLCELL_52_1295 ();
 FILLCELL_X32 FILLCELL_52_1327 ();
 FILLCELL_X32 FILLCELL_52_1359 ();
 FILLCELL_X32 FILLCELL_52_1391 ();
 FILLCELL_X32 FILLCELL_52_1423 ();
 FILLCELL_X32 FILLCELL_52_1455 ();
 FILLCELL_X32 FILLCELL_52_1487 ();
 FILLCELL_X32 FILLCELL_52_1519 ();
 FILLCELL_X32 FILLCELL_52_1551 ();
 FILLCELL_X32 FILLCELL_52_1583 ();
 FILLCELL_X32 FILLCELL_52_1615 ();
 FILLCELL_X32 FILLCELL_52_1647 ();
 FILLCELL_X32 FILLCELL_52_1679 ();
 FILLCELL_X32 FILLCELL_52_1711 ();
 FILLCELL_X32 FILLCELL_52_1743 ();
 FILLCELL_X32 FILLCELL_52_1775 ();
 FILLCELL_X32 FILLCELL_52_1807 ();
 FILLCELL_X32 FILLCELL_52_1839 ();
 FILLCELL_X16 FILLCELL_52_1871 ();
 FILLCELL_X8 FILLCELL_52_1887 ();
 FILLCELL_X2 FILLCELL_52_1895 ();
 FILLCELL_X32 FILLCELL_53_0 ();
 FILLCELL_X32 FILLCELL_53_32 ();
 FILLCELL_X32 FILLCELL_53_64 ();
 FILLCELL_X32 FILLCELL_53_96 ();
 FILLCELL_X32 FILLCELL_53_128 ();
 FILLCELL_X32 FILLCELL_53_160 ();
 FILLCELL_X32 FILLCELL_53_192 ();
 FILLCELL_X32 FILLCELL_53_224 ();
 FILLCELL_X32 FILLCELL_53_256 ();
 FILLCELL_X32 FILLCELL_53_288 ();
 FILLCELL_X32 FILLCELL_53_320 ();
 FILLCELL_X32 FILLCELL_53_352 ();
 FILLCELL_X32 FILLCELL_53_384 ();
 FILLCELL_X32 FILLCELL_53_416 ();
 FILLCELL_X32 FILLCELL_53_448 ();
 FILLCELL_X32 FILLCELL_53_480 ();
 FILLCELL_X16 FILLCELL_53_512 ();
 FILLCELL_X32 FILLCELL_53_532 ();
 FILLCELL_X32 FILLCELL_53_564 ();
 FILLCELL_X32 FILLCELL_53_596 ();
 FILLCELL_X32 FILLCELL_53_628 ();
 FILLCELL_X32 FILLCELL_53_660 ();
 FILLCELL_X32 FILLCELL_53_692 ();
 FILLCELL_X32 FILLCELL_53_724 ();
 FILLCELL_X32 FILLCELL_53_756 ();
 FILLCELL_X32 FILLCELL_53_788 ();
 FILLCELL_X32 FILLCELL_53_820 ();
 FILLCELL_X32 FILLCELL_53_852 ();
 FILLCELL_X32 FILLCELL_53_884 ();
 FILLCELL_X32 FILLCELL_53_916 ();
 FILLCELL_X32 FILLCELL_53_948 ();
 FILLCELL_X32 FILLCELL_53_980 ();
 FILLCELL_X32 FILLCELL_53_1012 ();
 FILLCELL_X32 FILLCELL_53_1044 ();
 FILLCELL_X32 FILLCELL_53_1076 ();
 FILLCELL_X32 FILLCELL_53_1108 ();
 FILLCELL_X32 FILLCELL_53_1140 ();
 FILLCELL_X32 FILLCELL_53_1172 ();
 FILLCELL_X32 FILLCELL_53_1204 ();
 FILLCELL_X32 FILLCELL_53_1236 ();
 FILLCELL_X32 FILLCELL_53_1268 ();
 FILLCELL_X32 FILLCELL_53_1300 ();
 FILLCELL_X32 FILLCELL_53_1332 ();
 FILLCELL_X32 FILLCELL_53_1364 ();
 FILLCELL_X32 FILLCELL_53_1396 ();
 FILLCELL_X32 FILLCELL_53_1428 ();
 FILLCELL_X32 FILLCELL_53_1460 ();
 FILLCELL_X32 FILLCELL_53_1492 ();
 FILLCELL_X32 FILLCELL_53_1524 ();
 FILLCELL_X32 FILLCELL_53_1556 ();
 FILLCELL_X32 FILLCELL_53_1588 ();
 FILLCELL_X32 FILLCELL_53_1620 ();
 FILLCELL_X32 FILLCELL_53_1652 ();
 FILLCELL_X32 FILLCELL_53_1684 ();
 FILLCELL_X32 FILLCELL_53_1716 ();
 FILLCELL_X32 FILLCELL_53_1748 ();
 FILLCELL_X32 FILLCELL_53_1780 ();
 FILLCELL_X32 FILLCELL_53_1812 ();
 FILLCELL_X32 FILLCELL_53_1844 ();
 FILLCELL_X16 FILLCELL_53_1876 ();
 FILLCELL_X4 FILLCELL_53_1892 ();
 FILLCELL_X1 FILLCELL_53_1896 ();
 FILLCELL_X32 FILLCELL_54_0 ();
 FILLCELL_X32 FILLCELL_54_32 ();
 FILLCELL_X32 FILLCELL_54_64 ();
 FILLCELL_X32 FILLCELL_54_96 ();
 FILLCELL_X32 FILLCELL_54_128 ();
 FILLCELL_X32 FILLCELL_54_160 ();
 FILLCELL_X32 FILLCELL_54_192 ();
 FILLCELL_X32 FILLCELL_54_224 ();
 FILLCELL_X32 FILLCELL_54_256 ();
 FILLCELL_X32 FILLCELL_54_288 ();
 FILLCELL_X32 FILLCELL_54_320 ();
 FILLCELL_X32 FILLCELL_54_352 ();
 FILLCELL_X32 FILLCELL_54_384 ();
 FILLCELL_X32 FILLCELL_54_416 ();
 FILLCELL_X32 FILLCELL_54_448 ();
 FILLCELL_X32 FILLCELL_54_483 ();
 FILLCELL_X32 FILLCELL_54_515 ();
 FILLCELL_X32 FILLCELL_54_547 ();
 FILLCELL_X32 FILLCELL_54_579 ();
 FILLCELL_X32 FILLCELL_54_611 ();
 FILLCELL_X32 FILLCELL_54_643 ();
 FILLCELL_X32 FILLCELL_54_675 ();
 FILLCELL_X32 FILLCELL_54_707 ();
 FILLCELL_X32 FILLCELL_54_739 ();
 FILLCELL_X32 FILLCELL_54_771 ();
 FILLCELL_X32 FILLCELL_54_803 ();
 FILLCELL_X32 FILLCELL_54_835 ();
 FILLCELL_X32 FILLCELL_54_867 ();
 FILLCELL_X32 FILLCELL_54_899 ();
 FILLCELL_X32 FILLCELL_54_931 ();
 FILLCELL_X32 FILLCELL_54_963 ();
 FILLCELL_X32 FILLCELL_54_995 ();
 FILLCELL_X32 FILLCELL_54_1027 ();
 FILLCELL_X32 FILLCELL_54_1059 ();
 FILLCELL_X32 FILLCELL_54_1091 ();
 FILLCELL_X32 FILLCELL_54_1123 ();
 FILLCELL_X32 FILLCELL_54_1155 ();
 FILLCELL_X32 FILLCELL_54_1187 ();
 FILLCELL_X32 FILLCELL_54_1219 ();
 FILLCELL_X32 FILLCELL_54_1251 ();
 FILLCELL_X32 FILLCELL_54_1283 ();
 FILLCELL_X32 FILLCELL_54_1315 ();
 FILLCELL_X32 FILLCELL_54_1347 ();
 FILLCELL_X32 FILLCELL_54_1379 ();
 FILLCELL_X32 FILLCELL_54_1411 ();
 FILLCELL_X32 FILLCELL_54_1443 ();
 FILLCELL_X32 FILLCELL_54_1475 ();
 FILLCELL_X32 FILLCELL_54_1507 ();
 FILLCELL_X32 FILLCELL_54_1539 ();
 FILLCELL_X32 FILLCELL_54_1571 ();
 FILLCELL_X32 FILLCELL_54_1603 ();
 FILLCELL_X32 FILLCELL_54_1635 ();
 FILLCELL_X32 FILLCELL_54_1667 ();
 FILLCELL_X32 FILLCELL_54_1699 ();
 FILLCELL_X32 FILLCELL_54_1731 ();
 FILLCELL_X32 FILLCELL_54_1763 ();
 FILLCELL_X32 FILLCELL_54_1795 ();
 FILLCELL_X32 FILLCELL_54_1827 ();
 FILLCELL_X32 FILLCELL_54_1859 ();
 FILLCELL_X4 FILLCELL_54_1891 ();
 FILLCELL_X2 FILLCELL_54_1895 ();
 FILLCELL_X32 FILLCELL_55_0 ();
 FILLCELL_X32 FILLCELL_55_32 ();
 FILLCELL_X32 FILLCELL_55_64 ();
 FILLCELL_X32 FILLCELL_55_96 ();
 FILLCELL_X32 FILLCELL_55_128 ();
 FILLCELL_X32 FILLCELL_55_160 ();
 FILLCELL_X32 FILLCELL_55_192 ();
 FILLCELL_X32 FILLCELL_55_224 ();
 FILLCELL_X32 FILLCELL_55_256 ();
 FILLCELL_X32 FILLCELL_55_288 ();
 FILLCELL_X32 FILLCELL_55_320 ();
 FILLCELL_X32 FILLCELL_55_352 ();
 FILLCELL_X32 FILLCELL_55_384 ();
 FILLCELL_X32 FILLCELL_55_416 ();
 FILLCELL_X32 FILLCELL_55_448 ();
 FILLCELL_X32 FILLCELL_55_480 ();
 FILLCELL_X8 FILLCELL_55_512 ();
 FILLCELL_X32 FILLCELL_55_524 ();
 FILLCELL_X32 FILLCELL_55_556 ();
 FILLCELL_X32 FILLCELL_55_588 ();
 FILLCELL_X32 FILLCELL_55_620 ();
 FILLCELL_X32 FILLCELL_55_652 ();
 FILLCELL_X4 FILLCELL_55_684 ();
 FILLCELL_X1 FILLCELL_55_688 ();
 FILLCELL_X32 FILLCELL_55_693 ();
 FILLCELL_X32 FILLCELL_55_725 ();
 FILLCELL_X32 FILLCELL_55_757 ();
 FILLCELL_X16 FILLCELL_55_789 ();
 FILLCELL_X4 FILLCELL_55_805 ();
 FILLCELL_X2 FILLCELL_55_809 ();
 FILLCELL_X1 FILLCELL_55_811 ();
 FILLCELL_X32 FILLCELL_55_816 ();
 FILLCELL_X32 FILLCELL_55_848 ();
 FILLCELL_X32 FILLCELL_55_880 ();
 FILLCELL_X32 FILLCELL_55_912 ();
 FILLCELL_X32 FILLCELL_55_944 ();
 FILLCELL_X32 FILLCELL_55_976 ();
 FILLCELL_X32 FILLCELL_55_1008 ();
 FILLCELL_X32 FILLCELL_55_1040 ();
 FILLCELL_X32 FILLCELL_55_1072 ();
 FILLCELL_X32 FILLCELL_55_1104 ();
 FILLCELL_X32 FILLCELL_55_1136 ();
 FILLCELL_X32 FILLCELL_55_1168 ();
 FILLCELL_X32 FILLCELL_55_1200 ();
 FILLCELL_X32 FILLCELL_55_1232 ();
 FILLCELL_X32 FILLCELL_55_1264 ();
 FILLCELL_X32 FILLCELL_55_1296 ();
 FILLCELL_X32 FILLCELL_55_1328 ();
 FILLCELL_X32 FILLCELL_55_1360 ();
 FILLCELL_X32 FILLCELL_55_1392 ();
 FILLCELL_X32 FILLCELL_55_1424 ();
 FILLCELL_X32 FILLCELL_55_1456 ();
 FILLCELL_X32 FILLCELL_55_1488 ();
 FILLCELL_X32 FILLCELL_55_1520 ();
 FILLCELL_X32 FILLCELL_55_1552 ();
 FILLCELL_X32 FILLCELL_55_1584 ();
 FILLCELL_X32 FILLCELL_55_1616 ();
 FILLCELL_X32 FILLCELL_55_1648 ();
 FILLCELL_X32 FILLCELL_55_1680 ();
 FILLCELL_X32 FILLCELL_55_1712 ();
 FILLCELL_X32 FILLCELL_55_1744 ();
 FILLCELL_X32 FILLCELL_55_1776 ();
 FILLCELL_X32 FILLCELL_55_1808 ();
 FILLCELL_X32 FILLCELL_55_1840 ();
 FILLCELL_X16 FILLCELL_55_1872 ();
 FILLCELL_X8 FILLCELL_55_1888 ();
 FILLCELL_X1 FILLCELL_55_1896 ();
 FILLCELL_X32 FILLCELL_56_0 ();
 FILLCELL_X32 FILLCELL_56_32 ();
 FILLCELL_X32 FILLCELL_56_64 ();
 FILLCELL_X32 FILLCELL_56_96 ();
 FILLCELL_X32 FILLCELL_56_128 ();
 FILLCELL_X32 FILLCELL_56_160 ();
 FILLCELL_X32 FILLCELL_56_192 ();
 FILLCELL_X32 FILLCELL_56_224 ();
 FILLCELL_X32 FILLCELL_56_256 ();
 FILLCELL_X32 FILLCELL_56_288 ();
 FILLCELL_X32 FILLCELL_56_320 ();
 FILLCELL_X32 FILLCELL_56_352 ();
 FILLCELL_X32 FILLCELL_56_384 ();
 FILLCELL_X32 FILLCELL_56_416 ();
 FILLCELL_X32 FILLCELL_56_448 ();
 FILLCELL_X32 FILLCELL_56_480 ();
 FILLCELL_X32 FILLCELL_56_512 ();
 FILLCELL_X32 FILLCELL_56_544 ();
 FILLCELL_X32 FILLCELL_56_576 ();
 FILLCELL_X32 FILLCELL_56_608 ();
 FILLCELL_X32 FILLCELL_56_640 ();
 FILLCELL_X16 FILLCELL_56_672 ();
 FILLCELL_X8 FILLCELL_56_688 ();
 FILLCELL_X4 FILLCELL_56_696 ();
 FILLCELL_X2 FILLCELL_56_700 ();
 FILLCELL_X4 FILLCELL_56_706 ();
 FILLCELL_X1 FILLCELL_56_710 ();
 FILLCELL_X32 FILLCELL_56_728 ();
 FILLCELL_X32 FILLCELL_56_760 ();
 FILLCELL_X16 FILLCELL_56_792 ();
 FILLCELL_X8 FILLCELL_56_808 ();
 FILLCELL_X4 FILLCELL_56_816 ();
 FILLCELL_X2 FILLCELL_56_820 ();
 FILLCELL_X8 FILLCELL_56_826 ();
 FILLCELL_X4 FILLCELL_56_834 ();
 FILLCELL_X2 FILLCELL_56_838 ();
 FILLCELL_X1 FILLCELL_56_840 ();
 FILLCELL_X32 FILLCELL_56_858 ();
 FILLCELL_X32 FILLCELL_56_890 ();
 FILLCELL_X32 FILLCELL_56_922 ();
 FILLCELL_X32 FILLCELL_56_954 ();
 FILLCELL_X32 FILLCELL_56_986 ();
 FILLCELL_X32 FILLCELL_56_1018 ();
 FILLCELL_X32 FILLCELL_56_1050 ();
 FILLCELL_X32 FILLCELL_56_1082 ();
 FILLCELL_X32 FILLCELL_56_1114 ();
 FILLCELL_X32 FILLCELL_56_1146 ();
 FILLCELL_X32 FILLCELL_56_1178 ();
 FILLCELL_X32 FILLCELL_56_1210 ();
 FILLCELL_X32 FILLCELL_56_1242 ();
 FILLCELL_X32 FILLCELL_56_1274 ();
 FILLCELL_X32 FILLCELL_56_1306 ();
 FILLCELL_X32 FILLCELL_56_1338 ();
 FILLCELL_X32 FILLCELL_56_1370 ();
 FILLCELL_X32 FILLCELL_56_1402 ();
 FILLCELL_X32 FILLCELL_56_1434 ();
 FILLCELL_X32 FILLCELL_56_1466 ();
 FILLCELL_X32 FILLCELL_56_1498 ();
 FILLCELL_X32 FILLCELL_56_1530 ();
 FILLCELL_X32 FILLCELL_56_1562 ();
 FILLCELL_X32 FILLCELL_56_1594 ();
 FILLCELL_X32 FILLCELL_56_1626 ();
 FILLCELL_X32 FILLCELL_56_1658 ();
 FILLCELL_X32 FILLCELL_56_1690 ();
 FILLCELL_X32 FILLCELL_56_1722 ();
 FILLCELL_X32 FILLCELL_56_1754 ();
 FILLCELL_X32 FILLCELL_56_1786 ();
 FILLCELL_X32 FILLCELL_56_1818 ();
 FILLCELL_X32 FILLCELL_56_1850 ();
 FILLCELL_X8 FILLCELL_56_1882 ();
 FILLCELL_X4 FILLCELL_56_1890 ();
 FILLCELL_X2 FILLCELL_56_1894 ();
 FILLCELL_X1 FILLCELL_56_1896 ();
 FILLCELL_X32 FILLCELL_57_0 ();
 FILLCELL_X32 FILLCELL_57_32 ();
 FILLCELL_X32 FILLCELL_57_64 ();
 FILLCELL_X32 FILLCELL_57_96 ();
 FILLCELL_X32 FILLCELL_57_128 ();
 FILLCELL_X32 FILLCELL_57_160 ();
 FILLCELL_X32 FILLCELL_57_192 ();
 FILLCELL_X32 FILLCELL_57_224 ();
 FILLCELL_X32 FILLCELL_57_256 ();
 FILLCELL_X32 FILLCELL_57_288 ();
 FILLCELL_X32 FILLCELL_57_320 ();
 FILLCELL_X32 FILLCELL_57_352 ();
 FILLCELL_X4 FILLCELL_57_384 ();
 FILLCELL_X32 FILLCELL_57_405 ();
 FILLCELL_X32 FILLCELL_57_437 ();
 FILLCELL_X32 FILLCELL_57_469 ();
 FILLCELL_X32 FILLCELL_57_501 ();
 FILLCELL_X32 FILLCELL_57_533 ();
 FILLCELL_X32 FILLCELL_57_565 ();
 FILLCELL_X32 FILLCELL_57_597 ();
 FILLCELL_X32 FILLCELL_57_629 ();
 FILLCELL_X16 FILLCELL_57_661 ();
 FILLCELL_X8 FILLCELL_57_677 ();
 FILLCELL_X1 FILLCELL_57_685 ();
 FILLCELL_X32 FILLCELL_57_689 ();
 FILLCELL_X32 FILLCELL_57_721 ();
 FILLCELL_X32 FILLCELL_57_753 ();
 FILLCELL_X32 FILLCELL_57_785 ();
 FILLCELL_X16 FILLCELL_57_817 ();
 FILLCELL_X4 FILLCELL_57_833 ();
 FILLCELL_X1 FILLCELL_57_837 ();
 FILLCELL_X32 FILLCELL_57_841 ();
 FILLCELL_X32 FILLCELL_57_873 ();
 FILLCELL_X32 FILLCELL_57_905 ();
 FILLCELL_X32 FILLCELL_57_937 ();
 FILLCELL_X32 FILLCELL_57_969 ();
 FILLCELL_X32 FILLCELL_57_1001 ();
 FILLCELL_X32 FILLCELL_57_1033 ();
 FILLCELL_X32 FILLCELL_57_1065 ();
 FILLCELL_X32 FILLCELL_57_1097 ();
 FILLCELL_X32 FILLCELL_57_1129 ();
 FILLCELL_X32 FILLCELL_57_1161 ();
 FILLCELL_X32 FILLCELL_57_1193 ();
 FILLCELL_X32 FILLCELL_57_1225 ();
 FILLCELL_X32 FILLCELL_57_1257 ();
 FILLCELL_X32 FILLCELL_57_1289 ();
 FILLCELL_X32 FILLCELL_57_1321 ();
 FILLCELL_X32 FILLCELL_57_1353 ();
 FILLCELL_X32 FILLCELL_57_1385 ();
 FILLCELL_X32 FILLCELL_57_1417 ();
 FILLCELL_X32 FILLCELL_57_1449 ();
 FILLCELL_X32 FILLCELL_57_1481 ();
 FILLCELL_X32 FILLCELL_57_1513 ();
 FILLCELL_X32 FILLCELL_57_1545 ();
 FILLCELL_X32 FILLCELL_57_1577 ();
 FILLCELL_X32 FILLCELL_57_1609 ();
 FILLCELL_X32 FILLCELL_57_1641 ();
 FILLCELL_X32 FILLCELL_57_1673 ();
 FILLCELL_X32 FILLCELL_57_1705 ();
 FILLCELL_X32 FILLCELL_57_1737 ();
 FILLCELL_X32 FILLCELL_57_1769 ();
 FILLCELL_X32 FILLCELL_57_1801 ();
 FILLCELL_X32 FILLCELL_57_1833 ();
 FILLCELL_X32 FILLCELL_57_1865 ();
 FILLCELL_X32 FILLCELL_58_0 ();
 FILLCELL_X32 FILLCELL_58_32 ();
 FILLCELL_X32 FILLCELL_58_64 ();
 FILLCELL_X32 FILLCELL_58_96 ();
 FILLCELL_X32 FILLCELL_58_128 ();
 FILLCELL_X32 FILLCELL_58_160 ();
 FILLCELL_X32 FILLCELL_58_192 ();
 FILLCELL_X32 FILLCELL_58_224 ();
 FILLCELL_X32 FILLCELL_58_256 ();
 FILLCELL_X32 FILLCELL_58_288 ();
 FILLCELL_X32 FILLCELL_58_320 ();
 FILLCELL_X32 FILLCELL_58_352 ();
 FILLCELL_X32 FILLCELL_58_384 ();
 FILLCELL_X32 FILLCELL_58_416 ();
 FILLCELL_X32 FILLCELL_58_448 ();
 FILLCELL_X32 FILLCELL_58_480 ();
 FILLCELL_X32 FILLCELL_58_512 ();
 FILLCELL_X32 FILLCELL_58_544 ();
 FILLCELL_X32 FILLCELL_58_576 ();
 FILLCELL_X32 FILLCELL_58_608 ();
 FILLCELL_X32 FILLCELL_58_640 ();
 FILLCELL_X32 FILLCELL_58_672 ();
 FILLCELL_X32 FILLCELL_58_704 ();
 FILLCELL_X32 FILLCELL_58_736 ();
 FILLCELL_X32 FILLCELL_58_768 ();
 FILLCELL_X32 FILLCELL_58_800 ();
 FILLCELL_X32 FILLCELL_58_832 ();
 FILLCELL_X32 FILLCELL_58_864 ();
 FILLCELL_X32 FILLCELL_58_896 ();
 FILLCELL_X32 FILLCELL_58_928 ();
 FILLCELL_X32 FILLCELL_58_960 ();
 FILLCELL_X32 FILLCELL_58_992 ();
 FILLCELL_X32 FILLCELL_58_1024 ();
 FILLCELL_X32 FILLCELL_58_1056 ();
 FILLCELL_X32 FILLCELL_58_1088 ();
 FILLCELL_X32 FILLCELL_58_1120 ();
 FILLCELL_X32 FILLCELL_58_1152 ();
 FILLCELL_X32 FILLCELL_58_1184 ();
 FILLCELL_X32 FILLCELL_58_1216 ();
 FILLCELL_X32 FILLCELL_58_1248 ();
 FILLCELL_X32 FILLCELL_58_1280 ();
 FILLCELL_X32 FILLCELL_58_1312 ();
 FILLCELL_X32 FILLCELL_58_1344 ();
 FILLCELL_X32 FILLCELL_58_1376 ();
 FILLCELL_X32 FILLCELL_58_1408 ();
 FILLCELL_X32 FILLCELL_58_1440 ();
 FILLCELL_X32 FILLCELL_58_1472 ();
 FILLCELL_X32 FILLCELL_58_1504 ();
 FILLCELL_X32 FILLCELL_58_1536 ();
 FILLCELL_X32 FILLCELL_58_1568 ();
 FILLCELL_X32 FILLCELL_58_1600 ();
 FILLCELL_X32 FILLCELL_58_1632 ();
 FILLCELL_X32 FILLCELL_58_1664 ();
 FILLCELL_X32 FILLCELL_58_1696 ();
 FILLCELL_X32 FILLCELL_58_1728 ();
 FILLCELL_X32 FILLCELL_58_1760 ();
 FILLCELL_X32 FILLCELL_58_1792 ();
 FILLCELL_X32 FILLCELL_58_1824 ();
 FILLCELL_X32 FILLCELL_58_1856 ();
 FILLCELL_X8 FILLCELL_58_1888 ();
 FILLCELL_X1 FILLCELL_58_1896 ();
 FILLCELL_X32 FILLCELL_59_0 ();
 FILLCELL_X32 FILLCELL_59_32 ();
 FILLCELL_X32 FILLCELL_59_64 ();
 FILLCELL_X32 FILLCELL_59_96 ();
 FILLCELL_X32 FILLCELL_59_128 ();
 FILLCELL_X32 FILLCELL_59_160 ();
 FILLCELL_X32 FILLCELL_59_192 ();
 FILLCELL_X32 FILLCELL_59_224 ();
 FILLCELL_X32 FILLCELL_59_256 ();
 FILLCELL_X32 FILLCELL_59_288 ();
 FILLCELL_X32 FILLCELL_59_320 ();
 FILLCELL_X32 FILLCELL_59_352 ();
 FILLCELL_X32 FILLCELL_59_384 ();
 FILLCELL_X32 FILLCELL_59_416 ();
 FILLCELL_X32 FILLCELL_59_448 ();
 FILLCELL_X32 FILLCELL_59_480 ();
 FILLCELL_X32 FILLCELL_59_512 ();
 FILLCELL_X32 FILLCELL_59_544 ();
 FILLCELL_X32 FILLCELL_59_576 ();
 FILLCELL_X32 FILLCELL_59_608 ();
 FILLCELL_X32 FILLCELL_59_640 ();
 FILLCELL_X32 FILLCELL_59_672 ();
 FILLCELL_X32 FILLCELL_59_704 ();
 FILLCELL_X32 FILLCELL_59_736 ();
 FILLCELL_X32 FILLCELL_59_768 ();
 FILLCELL_X32 FILLCELL_59_800 ();
 FILLCELL_X32 FILLCELL_59_832 ();
 FILLCELL_X32 FILLCELL_59_864 ();
 FILLCELL_X32 FILLCELL_59_896 ();
 FILLCELL_X32 FILLCELL_59_928 ();
 FILLCELL_X32 FILLCELL_59_960 ();
 FILLCELL_X32 FILLCELL_59_992 ();
 FILLCELL_X32 FILLCELL_59_1024 ();
 FILLCELL_X32 FILLCELL_59_1056 ();
 FILLCELL_X32 FILLCELL_59_1088 ();
 FILLCELL_X32 FILLCELL_59_1120 ();
 FILLCELL_X32 FILLCELL_59_1152 ();
 FILLCELL_X32 FILLCELL_59_1184 ();
 FILLCELL_X32 FILLCELL_59_1216 ();
 FILLCELL_X32 FILLCELL_59_1248 ();
 FILLCELL_X32 FILLCELL_59_1280 ();
 FILLCELL_X32 FILLCELL_59_1312 ();
 FILLCELL_X32 FILLCELL_59_1344 ();
 FILLCELL_X32 FILLCELL_59_1376 ();
 FILLCELL_X32 FILLCELL_59_1408 ();
 FILLCELL_X32 FILLCELL_59_1440 ();
 FILLCELL_X32 FILLCELL_59_1472 ();
 FILLCELL_X32 FILLCELL_59_1504 ();
 FILLCELL_X32 FILLCELL_59_1536 ();
 FILLCELL_X32 FILLCELL_59_1568 ();
 FILLCELL_X32 FILLCELL_59_1600 ();
 FILLCELL_X32 FILLCELL_59_1632 ();
 FILLCELL_X32 FILLCELL_59_1664 ();
 FILLCELL_X32 FILLCELL_59_1696 ();
 FILLCELL_X32 FILLCELL_59_1728 ();
 FILLCELL_X32 FILLCELL_59_1760 ();
 FILLCELL_X32 FILLCELL_59_1792 ();
 FILLCELL_X32 FILLCELL_59_1824 ();
 FILLCELL_X32 FILLCELL_59_1856 ();
 FILLCELL_X8 FILLCELL_59_1888 ();
 FILLCELL_X1 FILLCELL_59_1896 ();
 FILLCELL_X32 FILLCELL_60_0 ();
 FILLCELL_X32 FILLCELL_60_32 ();
 FILLCELL_X32 FILLCELL_60_64 ();
 FILLCELL_X32 FILLCELL_60_96 ();
 FILLCELL_X32 FILLCELL_60_128 ();
 FILLCELL_X32 FILLCELL_60_160 ();
 FILLCELL_X32 FILLCELL_60_192 ();
 FILLCELL_X32 FILLCELL_60_224 ();
 FILLCELL_X32 FILLCELL_60_256 ();
 FILLCELL_X32 FILLCELL_60_288 ();
 FILLCELL_X32 FILLCELL_60_320 ();
 FILLCELL_X32 FILLCELL_60_352 ();
 FILLCELL_X32 FILLCELL_60_384 ();
 FILLCELL_X32 FILLCELL_60_416 ();
 FILLCELL_X32 FILLCELL_60_448 ();
 FILLCELL_X32 FILLCELL_60_480 ();
 FILLCELL_X32 FILLCELL_60_512 ();
 FILLCELL_X32 FILLCELL_60_544 ();
 FILLCELL_X16 FILLCELL_60_576 ();
 FILLCELL_X8 FILLCELL_60_592 ();
 FILLCELL_X32 FILLCELL_60_617 ();
 FILLCELL_X32 FILLCELL_60_649 ();
 FILLCELL_X32 FILLCELL_60_681 ();
 FILLCELL_X32 FILLCELL_60_713 ();
 FILLCELL_X32 FILLCELL_60_745 ();
 FILLCELL_X32 FILLCELL_60_777 ();
 FILLCELL_X32 FILLCELL_60_809 ();
 FILLCELL_X32 FILLCELL_60_841 ();
 FILLCELL_X32 FILLCELL_60_873 ();
 FILLCELL_X32 FILLCELL_60_905 ();
 FILLCELL_X32 FILLCELL_60_937 ();
 FILLCELL_X32 FILLCELL_60_969 ();
 FILLCELL_X32 FILLCELL_60_1001 ();
 FILLCELL_X32 FILLCELL_60_1033 ();
 FILLCELL_X32 FILLCELL_60_1065 ();
 FILLCELL_X32 FILLCELL_60_1097 ();
 FILLCELL_X32 FILLCELL_60_1129 ();
 FILLCELL_X32 FILLCELL_60_1161 ();
 FILLCELL_X32 FILLCELL_60_1193 ();
 FILLCELL_X32 FILLCELL_60_1225 ();
 FILLCELL_X32 FILLCELL_60_1257 ();
 FILLCELL_X32 FILLCELL_60_1289 ();
 FILLCELL_X32 FILLCELL_60_1321 ();
 FILLCELL_X32 FILLCELL_60_1353 ();
 FILLCELL_X32 FILLCELL_60_1385 ();
 FILLCELL_X32 FILLCELL_60_1417 ();
 FILLCELL_X32 FILLCELL_60_1449 ();
 FILLCELL_X32 FILLCELL_60_1481 ();
 FILLCELL_X32 FILLCELL_60_1513 ();
 FILLCELL_X32 FILLCELL_60_1545 ();
 FILLCELL_X32 FILLCELL_60_1577 ();
 FILLCELL_X32 FILLCELL_60_1609 ();
 FILLCELL_X32 FILLCELL_60_1641 ();
 FILLCELL_X32 FILLCELL_60_1673 ();
 FILLCELL_X32 FILLCELL_60_1705 ();
 FILLCELL_X32 FILLCELL_60_1737 ();
 FILLCELL_X32 FILLCELL_60_1769 ();
 FILLCELL_X32 FILLCELL_60_1801 ();
 FILLCELL_X32 FILLCELL_60_1833 ();
 FILLCELL_X32 FILLCELL_60_1865 ();
 FILLCELL_X32 FILLCELL_61_0 ();
 FILLCELL_X32 FILLCELL_61_32 ();
 FILLCELL_X32 FILLCELL_61_64 ();
 FILLCELL_X32 FILLCELL_61_96 ();
 FILLCELL_X32 FILLCELL_61_128 ();
 FILLCELL_X32 FILLCELL_61_160 ();
 FILLCELL_X32 FILLCELL_61_192 ();
 FILLCELL_X32 FILLCELL_61_224 ();
 FILLCELL_X32 FILLCELL_61_256 ();
 FILLCELL_X16 FILLCELL_61_288 ();
 FILLCELL_X2 FILLCELL_61_304 ();
 FILLCELL_X32 FILLCELL_61_309 ();
 FILLCELL_X32 FILLCELL_61_341 ();
 FILLCELL_X32 FILLCELL_61_373 ();
 FILLCELL_X32 FILLCELL_61_405 ();
 FILLCELL_X32 FILLCELL_61_437 ();
 FILLCELL_X32 FILLCELL_61_469 ();
 FILLCELL_X32 FILLCELL_61_501 ();
 FILLCELL_X32 FILLCELL_61_533 ();
 FILLCELL_X32 FILLCELL_61_565 ();
 FILLCELL_X32 FILLCELL_61_597 ();
 FILLCELL_X32 FILLCELL_61_629 ();
 FILLCELL_X32 FILLCELL_61_661 ();
 FILLCELL_X32 FILLCELL_61_693 ();
 FILLCELL_X32 FILLCELL_61_725 ();
 FILLCELL_X32 FILLCELL_61_757 ();
 FILLCELL_X32 FILLCELL_61_789 ();
 FILLCELL_X32 FILLCELL_61_821 ();
 FILLCELL_X32 FILLCELL_61_853 ();
 FILLCELL_X32 FILLCELL_61_885 ();
 FILLCELL_X16 FILLCELL_61_917 ();
 FILLCELL_X4 FILLCELL_61_933 ();
 FILLCELL_X1 FILLCELL_61_937 ();
 FILLCELL_X32 FILLCELL_61_941 ();
 FILLCELL_X8 FILLCELL_61_973 ();
 FILLCELL_X32 FILLCELL_61_984 ();
 FILLCELL_X32 FILLCELL_61_1016 ();
 FILLCELL_X32 FILLCELL_61_1048 ();
 FILLCELL_X32 FILLCELL_61_1080 ();
 FILLCELL_X32 FILLCELL_61_1112 ();
 FILLCELL_X32 FILLCELL_61_1144 ();
 FILLCELL_X32 FILLCELL_61_1176 ();
 FILLCELL_X32 FILLCELL_61_1208 ();
 FILLCELL_X32 FILLCELL_61_1240 ();
 FILLCELL_X32 FILLCELL_61_1272 ();
 FILLCELL_X32 FILLCELL_61_1304 ();
 FILLCELL_X32 FILLCELL_61_1336 ();
 FILLCELL_X32 FILLCELL_61_1368 ();
 FILLCELL_X32 FILLCELL_61_1400 ();
 FILLCELL_X32 FILLCELL_61_1432 ();
 FILLCELL_X32 FILLCELL_61_1464 ();
 FILLCELL_X32 FILLCELL_61_1496 ();
 FILLCELL_X32 FILLCELL_61_1528 ();
 FILLCELL_X32 FILLCELL_61_1560 ();
 FILLCELL_X32 FILLCELL_61_1592 ();
 FILLCELL_X32 FILLCELL_61_1624 ();
 FILLCELL_X32 FILLCELL_61_1656 ();
 FILLCELL_X32 FILLCELL_61_1688 ();
 FILLCELL_X32 FILLCELL_61_1720 ();
 FILLCELL_X32 FILLCELL_61_1752 ();
 FILLCELL_X32 FILLCELL_61_1784 ();
 FILLCELL_X32 FILLCELL_61_1816 ();
 FILLCELL_X32 FILLCELL_61_1848 ();
 FILLCELL_X16 FILLCELL_61_1880 ();
 FILLCELL_X1 FILLCELL_61_1896 ();
 FILLCELL_X32 FILLCELL_62_0 ();
 FILLCELL_X32 FILLCELL_62_32 ();
 FILLCELL_X32 FILLCELL_62_64 ();
 FILLCELL_X32 FILLCELL_62_96 ();
 FILLCELL_X32 FILLCELL_62_128 ();
 FILLCELL_X32 FILLCELL_62_160 ();
 FILLCELL_X16 FILLCELL_62_192 ();
 FILLCELL_X4 FILLCELL_62_208 ();
 FILLCELL_X1 FILLCELL_62_212 ();
 FILLCELL_X32 FILLCELL_62_230 ();
 FILLCELL_X32 FILLCELL_62_262 ();
 FILLCELL_X32 FILLCELL_62_294 ();
 FILLCELL_X32 FILLCELL_62_326 ();
 FILLCELL_X32 FILLCELL_62_358 ();
 FILLCELL_X32 FILLCELL_62_390 ();
 FILLCELL_X32 FILLCELL_62_422 ();
 FILLCELL_X32 FILLCELL_62_454 ();
 FILLCELL_X32 FILLCELL_62_486 ();
 FILLCELL_X32 FILLCELL_62_518 ();
 FILLCELL_X32 FILLCELL_62_550 ();
 FILLCELL_X32 FILLCELL_62_582 ();
 FILLCELL_X32 FILLCELL_62_614 ();
 FILLCELL_X32 FILLCELL_62_646 ();
 FILLCELL_X32 FILLCELL_62_678 ();
 FILLCELL_X32 FILLCELL_62_710 ();
 FILLCELL_X32 FILLCELL_62_742 ();
 FILLCELL_X32 FILLCELL_62_774 ();
 FILLCELL_X32 FILLCELL_62_806 ();
 FILLCELL_X32 FILLCELL_62_838 ();
 FILLCELL_X32 FILLCELL_62_870 ();
 FILLCELL_X32 FILLCELL_62_902 ();
 FILLCELL_X32 FILLCELL_62_934 ();
 FILLCELL_X32 FILLCELL_62_966 ();
 FILLCELL_X32 FILLCELL_62_998 ();
 FILLCELL_X1 FILLCELL_62_1030 ();
 FILLCELL_X32 FILLCELL_62_1034 ();
 FILLCELL_X32 FILLCELL_62_1066 ();
 FILLCELL_X32 FILLCELL_62_1098 ();
 FILLCELL_X32 FILLCELL_62_1130 ();
 FILLCELL_X32 FILLCELL_62_1162 ();
 FILLCELL_X32 FILLCELL_62_1194 ();
 FILLCELL_X32 FILLCELL_62_1226 ();
 FILLCELL_X32 FILLCELL_62_1258 ();
 FILLCELL_X32 FILLCELL_62_1290 ();
 FILLCELL_X32 FILLCELL_62_1322 ();
 FILLCELL_X32 FILLCELL_62_1354 ();
 FILLCELL_X32 FILLCELL_62_1386 ();
 FILLCELL_X32 FILLCELL_62_1418 ();
 FILLCELL_X32 FILLCELL_62_1450 ();
 FILLCELL_X32 FILLCELL_62_1482 ();
 FILLCELL_X32 FILLCELL_62_1514 ();
 FILLCELL_X32 FILLCELL_62_1546 ();
 FILLCELL_X32 FILLCELL_62_1578 ();
 FILLCELL_X32 FILLCELL_62_1610 ();
 FILLCELL_X32 FILLCELL_62_1642 ();
 FILLCELL_X32 FILLCELL_62_1674 ();
 FILLCELL_X32 FILLCELL_62_1706 ();
 FILLCELL_X32 FILLCELL_62_1738 ();
 FILLCELL_X32 FILLCELL_62_1770 ();
 FILLCELL_X32 FILLCELL_62_1802 ();
 FILLCELL_X32 FILLCELL_62_1834 ();
 FILLCELL_X16 FILLCELL_62_1866 ();
 FILLCELL_X8 FILLCELL_62_1882 ();
 FILLCELL_X4 FILLCELL_62_1890 ();
 FILLCELL_X2 FILLCELL_62_1894 ();
 FILLCELL_X1 FILLCELL_62_1896 ();
 FILLCELL_X32 FILLCELL_63_0 ();
 FILLCELL_X32 FILLCELL_63_32 ();
 FILLCELL_X32 FILLCELL_63_64 ();
 FILLCELL_X32 FILLCELL_63_96 ();
 FILLCELL_X32 FILLCELL_63_128 ();
 FILLCELL_X32 FILLCELL_63_160 ();
 FILLCELL_X32 FILLCELL_63_192 ();
 FILLCELL_X32 FILLCELL_63_224 ();
 FILLCELL_X32 FILLCELL_63_256 ();
 FILLCELL_X32 FILLCELL_63_288 ();
 FILLCELL_X32 FILLCELL_63_320 ();
 FILLCELL_X32 FILLCELL_63_352 ();
 FILLCELL_X32 FILLCELL_63_384 ();
 FILLCELL_X32 FILLCELL_63_416 ();
 FILLCELL_X32 FILLCELL_63_448 ();
 FILLCELL_X32 FILLCELL_63_480 ();
 FILLCELL_X32 FILLCELL_63_512 ();
 FILLCELL_X32 FILLCELL_63_544 ();
 FILLCELL_X32 FILLCELL_63_576 ();
 FILLCELL_X32 FILLCELL_63_608 ();
 FILLCELL_X32 FILLCELL_63_640 ();
 FILLCELL_X32 FILLCELL_63_672 ();
 FILLCELL_X32 FILLCELL_63_704 ();
 FILLCELL_X32 FILLCELL_63_736 ();
 FILLCELL_X32 FILLCELL_63_768 ();
 FILLCELL_X32 FILLCELL_63_800 ();
 FILLCELL_X32 FILLCELL_63_832 ();
 FILLCELL_X32 FILLCELL_63_864 ();
 FILLCELL_X32 FILLCELL_63_896 ();
 FILLCELL_X32 FILLCELL_63_928 ();
 FILLCELL_X32 FILLCELL_63_960 ();
 FILLCELL_X32 FILLCELL_63_992 ();
 FILLCELL_X32 FILLCELL_63_1024 ();
 FILLCELL_X8 FILLCELL_63_1056 ();
 FILLCELL_X2 FILLCELL_63_1064 ();
 FILLCELL_X1 FILLCELL_63_1066 ();
 FILLCELL_X32 FILLCELL_63_1070 ();
 FILLCELL_X32 FILLCELL_63_1102 ();
 FILLCELL_X32 FILLCELL_63_1134 ();
 FILLCELL_X32 FILLCELL_63_1166 ();
 FILLCELL_X32 FILLCELL_63_1198 ();
 FILLCELL_X32 FILLCELL_63_1230 ();
 FILLCELL_X32 FILLCELL_63_1262 ();
 FILLCELL_X32 FILLCELL_63_1294 ();
 FILLCELL_X32 FILLCELL_63_1326 ();
 FILLCELL_X32 FILLCELL_63_1358 ();
 FILLCELL_X32 FILLCELL_63_1390 ();
 FILLCELL_X32 FILLCELL_63_1422 ();
 FILLCELL_X32 FILLCELL_63_1454 ();
 FILLCELL_X32 FILLCELL_63_1486 ();
 FILLCELL_X32 FILLCELL_63_1518 ();
 FILLCELL_X32 FILLCELL_63_1550 ();
 FILLCELL_X32 FILLCELL_63_1582 ();
 FILLCELL_X32 FILLCELL_63_1614 ();
 FILLCELL_X32 FILLCELL_63_1646 ();
 FILLCELL_X32 FILLCELL_63_1678 ();
 FILLCELL_X32 FILLCELL_63_1710 ();
 FILLCELL_X32 FILLCELL_63_1742 ();
 FILLCELL_X32 FILLCELL_63_1774 ();
 FILLCELL_X32 FILLCELL_63_1806 ();
 FILLCELL_X32 FILLCELL_63_1838 ();
 FILLCELL_X16 FILLCELL_63_1870 ();
 FILLCELL_X8 FILLCELL_63_1886 ();
 FILLCELL_X2 FILLCELL_63_1894 ();
 FILLCELL_X1 FILLCELL_63_1896 ();
 FILLCELL_X32 FILLCELL_64_0 ();
 FILLCELL_X32 FILLCELL_64_32 ();
 FILLCELL_X32 FILLCELL_64_64 ();
 FILLCELL_X32 FILLCELL_64_96 ();
 FILLCELL_X32 FILLCELL_64_128 ();
 FILLCELL_X32 FILLCELL_64_160 ();
 FILLCELL_X32 FILLCELL_64_192 ();
 FILLCELL_X32 FILLCELL_64_224 ();
 FILLCELL_X16 FILLCELL_64_256 ();
 FILLCELL_X8 FILLCELL_64_272 ();
 FILLCELL_X2 FILLCELL_64_280 ();
 FILLCELL_X1 FILLCELL_64_282 ();
 FILLCELL_X32 FILLCELL_64_290 ();
 FILLCELL_X32 FILLCELL_64_322 ();
 FILLCELL_X32 FILLCELL_64_354 ();
 FILLCELL_X32 FILLCELL_64_386 ();
 FILLCELL_X32 FILLCELL_64_418 ();
 FILLCELL_X32 FILLCELL_64_450 ();
 FILLCELL_X32 FILLCELL_64_482 ();
 FILLCELL_X32 FILLCELL_64_514 ();
 FILLCELL_X32 FILLCELL_64_546 ();
 FILLCELL_X32 FILLCELL_64_578 ();
 FILLCELL_X32 FILLCELL_64_610 ();
 FILLCELL_X32 FILLCELL_64_642 ();
 FILLCELL_X32 FILLCELL_64_674 ();
 FILLCELL_X32 FILLCELL_64_706 ();
 FILLCELL_X32 FILLCELL_64_738 ();
 FILLCELL_X32 FILLCELL_64_770 ();
 FILLCELL_X32 FILLCELL_64_802 ();
 FILLCELL_X32 FILLCELL_64_834 ();
 FILLCELL_X32 FILLCELL_64_866 ();
 FILLCELL_X32 FILLCELL_64_898 ();
 FILLCELL_X32 FILLCELL_64_930 ();
 FILLCELL_X32 FILLCELL_64_962 ();
 FILLCELL_X32 FILLCELL_64_994 ();
 FILLCELL_X32 FILLCELL_64_1026 ();
 FILLCELL_X32 FILLCELL_64_1058 ();
 FILLCELL_X32 FILLCELL_64_1090 ();
 FILLCELL_X32 FILLCELL_64_1122 ();
 FILLCELL_X32 FILLCELL_64_1154 ();
 FILLCELL_X32 FILLCELL_64_1186 ();
 FILLCELL_X32 FILLCELL_64_1218 ();
 FILLCELL_X32 FILLCELL_64_1250 ();
 FILLCELL_X32 FILLCELL_64_1282 ();
 FILLCELL_X32 FILLCELL_64_1314 ();
 FILLCELL_X32 FILLCELL_64_1346 ();
 FILLCELL_X32 FILLCELL_64_1378 ();
 FILLCELL_X32 FILLCELL_64_1410 ();
 FILLCELL_X32 FILLCELL_64_1442 ();
 FILLCELL_X32 FILLCELL_64_1474 ();
 FILLCELL_X32 FILLCELL_64_1506 ();
 FILLCELL_X32 FILLCELL_64_1538 ();
 FILLCELL_X32 FILLCELL_64_1570 ();
 FILLCELL_X32 FILLCELL_64_1602 ();
 FILLCELL_X32 FILLCELL_64_1634 ();
 FILLCELL_X32 FILLCELL_64_1666 ();
 FILLCELL_X32 FILLCELL_64_1698 ();
 FILLCELL_X32 FILLCELL_64_1730 ();
 FILLCELL_X32 FILLCELL_64_1762 ();
 FILLCELL_X32 FILLCELL_64_1794 ();
 FILLCELL_X32 FILLCELL_64_1826 ();
 FILLCELL_X32 FILLCELL_64_1858 ();
 FILLCELL_X4 FILLCELL_64_1890 ();
 FILLCELL_X2 FILLCELL_64_1894 ();
 FILLCELL_X1 FILLCELL_64_1896 ();
 FILLCELL_X32 FILLCELL_65_0 ();
 FILLCELL_X32 FILLCELL_65_32 ();
 FILLCELL_X32 FILLCELL_65_64 ();
 FILLCELL_X32 FILLCELL_65_96 ();
 FILLCELL_X32 FILLCELL_65_128 ();
 FILLCELL_X32 FILLCELL_65_160 ();
 FILLCELL_X32 FILLCELL_65_192 ();
 FILLCELL_X32 FILLCELL_65_224 ();
 FILLCELL_X32 FILLCELL_65_256 ();
 FILLCELL_X2 FILLCELL_65_288 ();
 FILLCELL_X1 FILLCELL_65_290 ();
 FILLCELL_X2 FILLCELL_65_294 ();
 FILLCELL_X32 FILLCELL_65_301 ();
 FILLCELL_X32 FILLCELL_65_333 ();
 FILLCELL_X32 FILLCELL_65_365 ();
 FILLCELL_X8 FILLCELL_65_397 ();
 FILLCELL_X32 FILLCELL_65_412 ();
 FILLCELL_X32 FILLCELL_65_444 ();
 FILLCELL_X32 FILLCELL_65_476 ();
 FILLCELL_X32 FILLCELL_65_508 ();
 FILLCELL_X32 FILLCELL_65_540 ();
 FILLCELL_X32 FILLCELL_65_572 ();
 FILLCELL_X8 FILLCELL_65_604 ();
 FILLCELL_X2 FILLCELL_65_612 ();
 FILLCELL_X1 FILLCELL_65_614 ();
 FILLCELL_X32 FILLCELL_65_622 ();
 FILLCELL_X32 FILLCELL_65_654 ();
 FILLCELL_X32 FILLCELL_65_686 ();
 FILLCELL_X32 FILLCELL_65_718 ();
 FILLCELL_X32 FILLCELL_65_750 ();
 FILLCELL_X32 FILLCELL_65_782 ();
 FILLCELL_X32 FILLCELL_65_814 ();
 FILLCELL_X32 FILLCELL_65_846 ();
 FILLCELL_X8 FILLCELL_65_878 ();
 FILLCELL_X4 FILLCELL_65_886 ();
 FILLCELL_X2 FILLCELL_65_890 ();
 FILLCELL_X32 FILLCELL_65_895 ();
 FILLCELL_X32 FILLCELL_65_927 ();
 FILLCELL_X32 FILLCELL_65_959 ();
 FILLCELL_X32 FILLCELL_65_991 ();
 FILLCELL_X32 FILLCELL_65_1023 ();
 FILLCELL_X32 FILLCELL_65_1055 ();
 FILLCELL_X32 FILLCELL_65_1087 ();
 FILLCELL_X32 FILLCELL_65_1119 ();
 FILLCELL_X32 FILLCELL_65_1151 ();
 FILLCELL_X32 FILLCELL_65_1183 ();
 FILLCELL_X32 FILLCELL_65_1215 ();
 FILLCELL_X32 FILLCELL_65_1247 ();
 FILLCELL_X32 FILLCELL_65_1279 ();
 FILLCELL_X32 FILLCELL_65_1311 ();
 FILLCELL_X32 FILLCELL_65_1343 ();
 FILLCELL_X32 FILLCELL_65_1375 ();
 FILLCELL_X32 FILLCELL_65_1407 ();
 FILLCELL_X32 FILLCELL_65_1439 ();
 FILLCELL_X32 FILLCELL_65_1471 ();
 FILLCELL_X32 FILLCELL_65_1503 ();
 FILLCELL_X32 FILLCELL_65_1535 ();
 FILLCELL_X32 FILLCELL_65_1567 ();
 FILLCELL_X32 FILLCELL_65_1599 ();
 FILLCELL_X32 FILLCELL_65_1631 ();
 FILLCELL_X32 FILLCELL_65_1663 ();
 FILLCELL_X32 FILLCELL_65_1695 ();
 FILLCELL_X32 FILLCELL_65_1727 ();
 FILLCELL_X32 FILLCELL_65_1759 ();
 FILLCELL_X32 FILLCELL_65_1791 ();
 FILLCELL_X32 FILLCELL_65_1823 ();
 FILLCELL_X32 FILLCELL_65_1855 ();
 FILLCELL_X8 FILLCELL_65_1887 ();
 FILLCELL_X2 FILLCELL_65_1895 ();
 FILLCELL_X32 FILLCELL_66_0 ();
 FILLCELL_X32 FILLCELL_66_32 ();
 FILLCELL_X32 FILLCELL_66_64 ();
 FILLCELL_X32 FILLCELL_66_96 ();
 FILLCELL_X32 FILLCELL_66_128 ();
 FILLCELL_X32 FILLCELL_66_160 ();
 FILLCELL_X32 FILLCELL_66_192 ();
 FILLCELL_X32 FILLCELL_66_224 ();
 FILLCELL_X32 FILLCELL_66_256 ();
 FILLCELL_X16 FILLCELL_66_288 ();
 FILLCELL_X4 FILLCELL_66_304 ();
 FILLCELL_X2 FILLCELL_66_308 ();
 FILLCELL_X32 FILLCELL_66_314 ();
 FILLCELL_X32 FILLCELL_66_346 ();
 FILLCELL_X32 FILLCELL_66_378 ();
 FILLCELL_X32 FILLCELL_66_410 ();
 FILLCELL_X32 FILLCELL_66_442 ();
 FILLCELL_X32 FILLCELL_66_474 ();
 FILLCELL_X32 FILLCELL_66_506 ();
 FILLCELL_X32 FILLCELL_66_538 ();
 FILLCELL_X32 FILLCELL_66_570 ();
 FILLCELL_X32 FILLCELL_66_602 ();
 FILLCELL_X32 FILLCELL_66_634 ();
 FILLCELL_X32 FILLCELL_66_666 ();
 FILLCELL_X32 FILLCELL_66_698 ();
 FILLCELL_X32 FILLCELL_66_730 ();
 FILLCELL_X32 FILLCELL_66_762 ();
 FILLCELL_X32 FILLCELL_66_794 ();
 FILLCELL_X32 FILLCELL_66_826 ();
 FILLCELL_X32 FILLCELL_66_858 ();
 FILLCELL_X32 FILLCELL_66_890 ();
 FILLCELL_X32 FILLCELL_66_922 ();
 FILLCELL_X32 FILLCELL_66_954 ();
 FILLCELL_X32 FILLCELL_66_986 ();
 FILLCELL_X4 FILLCELL_66_1018 ();
 FILLCELL_X32 FILLCELL_66_1027 ();
 FILLCELL_X32 FILLCELL_66_1059 ();
 FILLCELL_X32 FILLCELL_66_1091 ();
 FILLCELL_X32 FILLCELL_66_1123 ();
 FILLCELL_X32 FILLCELL_66_1155 ();
 FILLCELL_X32 FILLCELL_66_1187 ();
 FILLCELL_X32 FILLCELL_66_1219 ();
 FILLCELL_X32 FILLCELL_66_1251 ();
 FILLCELL_X32 FILLCELL_66_1283 ();
 FILLCELL_X32 FILLCELL_66_1315 ();
 FILLCELL_X32 FILLCELL_66_1347 ();
 FILLCELL_X32 FILLCELL_66_1379 ();
 FILLCELL_X32 FILLCELL_66_1411 ();
 FILLCELL_X32 FILLCELL_66_1443 ();
 FILLCELL_X32 FILLCELL_66_1475 ();
 FILLCELL_X32 FILLCELL_66_1507 ();
 FILLCELL_X32 FILLCELL_66_1539 ();
 FILLCELL_X32 FILLCELL_66_1571 ();
 FILLCELL_X32 FILLCELL_66_1603 ();
 FILLCELL_X32 FILLCELL_66_1635 ();
 FILLCELL_X32 FILLCELL_66_1667 ();
 FILLCELL_X32 FILLCELL_66_1699 ();
 FILLCELL_X32 FILLCELL_66_1731 ();
 FILLCELL_X32 FILLCELL_66_1763 ();
 FILLCELL_X32 FILLCELL_66_1795 ();
 FILLCELL_X32 FILLCELL_66_1827 ();
 FILLCELL_X32 FILLCELL_66_1859 ();
 FILLCELL_X4 FILLCELL_66_1891 ();
 FILLCELL_X2 FILLCELL_66_1895 ();
 FILLCELL_X32 FILLCELL_67_0 ();
 FILLCELL_X32 FILLCELL_67_32 ();
 FILLCELL_X32 FILLCELL_67_64 ();
 FILLCELL_X32 FILLCELL_67_96 ();
 FILLCELL_X32 FILLCELL_67_128 ();
 FILLCELL_X32 FILLCELL_67_160 ();
 FILLCELL_X32 FILLCELL_67_192 ();
 FILLCELL_X32 FILLCELL_67_224 ();
 FILLCELL_X32 FILLCELL_67_256 ();
 FILLCELL_X32 FILLCELL_67_288 ();
 FILLCELL_X32 FILLCELL_67_320 ();
 FILLCELL_X32 FILLCELL_67_352 ();
 FILLCELL_X16 FILLCELL_67_384 ();
 FILLCELL_X8 FILLCELL_67_400 ();
 FILLCELL_X4 FILLCELL_67_408 ();
 FILLCELL_X2 FILLCELL_67_412 ();
 FILLCELL_X1 FILLCELL_67_414 ();
 FILLCELL_X32 FILLCELL_67_418 ();
 FILLCELL_X32 FILLCELL_67_450 ();
 FILLCELL_X16 FILLCELL_67_482 ();
 FILLCELL_X2 FILLCELL_67_498 ();
 FILLCELL_X32 FILLCELL_67_502 ();
 FILLCELL_X32 FILLCELL_67_534 ();
 FILLCELL_X32 FILLCELL_67_566 ();
 FILLCELL_X4 FILLCELL_67_598 ();
 FILLCELL_X32 FILLCELL_67_604 ();
 FILLCELL_X32 FILLCELL_67_636 ();
 FILLCELL_X32 FILLCELL_67_668 ();
 FILLCELL_X32 FILLCELL_67_700 ();
 FILLCELL_X32 FILLCELL_67_732 ();
 FILLCELL_X32 FILLCELL_67_764 ();
 FILLCELL_X32 FILLCELL_67_796 ();
 FILLCELL_X32 FILLCELL_67_828 ();
 FILLCELL_X32 FILLCELL_67_860 ();
 FILLCELL_X32 FILLCELL_67_892 ();
 FILLCELL_X32 FILLCELL_67_924 ();
 FILLCELL_X32 FILLCELL_67_956 ();
 FILLCELL_X32 FILLCELL_67_988 ();
 FILLCELL_X16 FILLCELL_67_1020 ();
 FILLCELL_X2 FILLCELL_67_1036 ();
 FILLCELL_X1 FILLCELL_67_1038 ();
 FILLCELL_X32 FILLCELL_67_1043 ();
 FILLCELL_X32 FILLCELL_67_1075 ();
 FILLCELL_X32 FILLCELL_67_1107 ();
 FILLCELL_X32 FILLCELL_67_1139 ();
 FILLCELL_X32 FILLCELL_67_1171 ();
 FILLCELL_X32 FILLCELL_67_1203 ();
 FILLCELL_X32 FILLCELL_67_1235 ();
 FILLCELL_X32 FILLCELL_67_1267 ();
 FILLCELL_X32 FILLCELL_67_1299 ();
 FILLCELL_X32 FILLCELL_67_1331 ();
 FILLCELL_X32 FILLCELL_67_1363 ();
 FILLCELL_X32 FILLCELL_67_1395 ();
 FILLCELL_X32 FILLCELL_67_1427 ();
 FILLCELL_X32 FILLCELL_67_1459 ();
 FILLCELL_X32 FILLCELL_67_1491 ();
 FILLCELL_X32 FILLCELL_67_1523 ();
 FILLCELL_X32 FILLCELL_67_1555 ();
 FILLCELL_X32 FILLCELL_67_1587 ();
 FILLCELL_X32 FILLCELL_67_1619 ();
 FILLCELL_X32 FILLCELL_67_1651 ();
 FILLCELL_X32 FILLCELL_67_1683 ();
 FILLCELL_X32 FILLCELL_67_1715 ();
 FILLCELL_X32 FILLCELL_67_1747 ();
 FILLCELL_X32 FILLCELL_67_1779 ();
 FILLCELL_X32 FILLCELL_67_1811 ();
 FILLCELL_X32 FILLCELL_67_1843 ();
 FILLCELL_X16 FILLCELL_67_1875 ();
 FILLCELL_X4 FILLCELL_67_1891 ();
 FILLCELL_X2 FILLCELL_67_1895 ();
 FILLCELL_X32 FILLCELL_68_0 ();
 FILLCELL_X32 FILLCELL_68_32 ();
 FILLCELL_X32 FILLCELL_68_64 ();
 FILLCELL_X32 FILLCELL_68_96 ();
 FILLCELL_X32 FILLCELL_68_128 ();
 FILLCELL_X32 FILLCELL_68_160 ();
 FILLCELL_X32 FILLCELL_68_192 ();
 FILLCELL_X32 FILLCELL_68_224 ();
 FILLCELL_X32 FILLCELL_68_256 ();
 FILLCELL_X32 FILLCELL_68_288 ();
 FILLCELL_X32 FILLCELL_68_320 ();
 FILLCELL_X32 FILLCELL_68_352 ();
 FILLCELL_X32 FILLCELL_68_384 ();
 FILLCELL_X32 FILLCELL_68_416 ();
 FILLCELL_X16 FILLCELL_68_448 ();
 FILLCELL_X4 FILLCELL_68_464 ();
 FILLCELL_X1 FILLCELL_68_468 ();
 FILLCELL_X8 FILLCELL_68_474 ();
 FILLCELL_X2 FILLCELL_68_482 ();
 FILLCELL_X1 FILLCELL_68_484 ();
 FILLCELL_X32 FILLCELL_68_490 ();
 FILLCELL_X32 FILLCELL_68_522 ();
 FILLCELL_X32 FILLCELL_68_554 ();
 FILLCELL_X32 FILLCELL_68_586 ();
 FILLCELL_X32 FILLCELL_68_618 ();
 FILLCELL_X32 FILLCELL_68_650 ();
 FILLCELL_X32 FILLCELL_68_682 ();
 FILLCELL_X32 FILLCELL_68_714 ();
 FILLCELL_X32 FILLCELL_68_746 ();
 FILLCELL_X32 FILLCELL_68_778 ();
 FILLCELL_X32 FILLCELL_68_810 ();
 FILLCELL_X32 FILLCELL_68_842 ();
 FILLCELL_X32 FILLCELL_68_874 ();
 FILLCELL_X32 FILLCELL_68_906 ();
 FILLCELL_X32 FILLCELL_68_938 ();
 FILLCELL_X32 FILLCELL_68_970 ();
 FILLCELL_X32 FILLCELL_68_1002 ();
 FILLCELL_X32 FILLCELL_68_1034 ();
 FILLCELL_X32 FILLCELL_68_1066 ();
 FILLCELL_X32 FILLCELL_68_1098 ();
 FILLCELL_X32 FILLCELL_68_1130 ();
 FILLCELL_X32 FILLCELL_68_1162 ();
 FILLCELL_X32 FILLCELL_68_1194 ();
 FILLCELL_X32 FILLCELL_68_1226 ();
 FILLCELL_X32 FILLCELL_68_1258 ();
 FILLCELL_X32 FILLCELL_68_1290 ();
 FILLCELL_X32 FILLCELL_68_1322 ();
 FILLCELL_X32 FILLCELL_68_1354 ();
 FILLCELL_X32 FILLCELL_68_1386 ();
 FILLCELL_X32 FILLCELL_68_1418 ();
 FILLCELL_X32 FILLCELL_68_1450 ();
 FILLCELL_X32 FILLCELL_68_1482 ();
 FILLCELL_X32 FILLCELL_68_1514 ();
 FILLCELL_X32 FILLCELL_68_1546 ();
 FILLCELL_X32 FILLCELL_68_1578 ();
 FILLCELL_X32 FILLCELL_68_1610 ();
 FILLCELL_X32 FILLCELL_68_1642 ();
 FILLCELL_X32 FILLCELL_68_1674 ();
 FILLCELL_X32 FILLCELL_68_1706 ();
 FILLCELL_X32 FILLCELL_68_1738 ();
 FILLCELL_X32 FILLCELL_68_1770 ();
 FILLCELL_X32 FILLCELL_68_1802 ();
 FILLCELL_X32 FILLCELL_68_1834 ();
 FILLCELL_X16 FILLCELL_68_1866 ();
 FILLCELL_X8 FILLCELL_68_1882 ();
 FILLCELL_X4 FILLCELL_68_1890 ();
 FILLCELL_X2 FILLCELL_68_1894 ();
 FILLCELL_X1 FILLCELL_68_1896 ();
 FILLCELL_X32 FILLCELL_69_0 ();
 FILLCELL_X32 FILLCELL_69_32 ();
 FILLCELL_X32 FILLCELL_69_64 ();
 FILLCELL_X32 FILLCELL_69_96 ();
 FILLCELL_X32 FILLCELL_69_128 ();
 FILLCELL_X32 FILLCELL_69_160 ();
 FILLCELL_X32 FILLCELL_69_192 ();
 FILLCELL_X32 FILLCELL_69_224 ();
 FILLCELL_X32 FILLCELL_69_256 ();
 FILLCELL_X32 FILLCELL_69_288 ();
 FILLCELL_X32 FILLCELL_69_320 ();
 FILLCELL_X32 FILLCELL_69_352 ();
 FILLCELL_X32 FILLCELL_69_384 ();
 FILLCELL_X32 FILLCELL_69_416 ();
 FILLCELL_X32 FILLCELL_69_448 ();
 FILLCELL_X32 FILLCELL_69_480 ();
 FILLCELL_X32 FILLCELL_69_516 ();
 FILLCELL_X32 FILLCELL_69_548 ();
 FILLCELL_X32 FILLCELL_69_580 ();
 FILLCELL_X32 FILLCELL_69_612 ();
 FILLCELL_X32 FILLCELL_69_644 ();
 FILLCELL_X32 FILLCELL_69_676 ();
 FILLCELL_X32 FILLCELL_69_708 ();
 FILLCELL_X32 FILLCELL_69_740 ();
 FILLCELL_X32 FILLCELL_69_772 ();
 FILLCELL_X32 FILLCELL_69_804 ();
 FILLCELL_X32 FILLCELL_69_836 ();
 FILLCELL_X32 FILLCELL_69_868 ();
 FILLCELL_X32 FILLCELL_69_900 ();
 FILLCELL_X32 FILLCELL_69_932 ();
 FILLCELL_X32 FILLCELL_69_964 ();
 FILLCELL_X32 FILLCELL_69_996 ();
 FILLCELL_X32 FILLCELL_69_1028 ();
 FILLCELL_X32 FILLCELL_69_1060 ();
 FILLCELL_X32 FILLCELL_69_1092 ();
 FILLCELL_X32 FILLCELL_69_1124 ();
 FILLCELL_X32 FILLCELL_69_1156 ();
 FILLCELL_X32 FILLCELL_69_1188 ();
 FILLCELL_X32 FILLCELL_69_1220 ();
 FILLCELL_X32 FILLCELL_69_1252 ();
 FILLCELL_X32 FILLCELL_69_1284 ();
 FILLCELL_X32 FILLCELL_69_1316 ();
 FILLCELL_X32 FILLCELL_69_1348 ();
 FILLCELL_X32 FILLCELL_69_1380 ();
 FILLCELL_X32 FILLCELL_69_1412 ();
 FILLCELL_X32 FILLCELL_69_1444 ();
 FILLCELL_X32 FILLCELL_69_1476 ();
 FILLCELL_X32 FILLCELL_69_1508 ();
 FILLCELL_X32 FILLCELL_69_1540 ();
 FILLCELL_X32 FILLCELL_69_1572 ();
 FILLCELL_X32 FILLCELL_69_1604 ();
 FILLCELL_X32 FILLCELL_69_1636 ();
 FILLCELL_X32 FILLCELL_69_1668 ();
 FILLCELL_X32 FILLCELL_69_1700 ();
 FILLCELL_X32 FILLCELL_69_1732 ();
 FILLCELL_X32 FILLCELL_69_1764 ();
 FILLCELL_X32 FILLCELL_69_1796 ();
 FILLCELL_X32 FILLCELL_69_1828 ();
 FILLCELL_X32 FILLCELL_69_1860 ();
 FILLCELL_X4 FILLCELL_69_1892 ();
 FILLCELL_X1 FILLCELL_69_1896 ();
 FILLCELL_X32 FILLCELL_70_0 ();
 FILLCELL_X32 FILLCELL_70_32 ();
 FILLCELL_X32 FILLCELL_70_64 ();
 FILLCELL_X32 FILLCELL_70_96 ();
 FILLCELL_X32 FILLCELL_70_128 ();
 FILLCELL_X32 FILLCELL_70_160 ();
 FILLCELL_X32 FILLCELL_70_192 ();
 FILLCELL_X32 FILLCELL_70_224 ();
 FILLCELL_X32 FILLCELL_70_256 ();
 FILLCELL_X32 FILLCELL_70_288 ();
 FILLCELL_X32 FILLCELL_70_320 ();
 FILLCELL_X32 FILLCELL_70_352 ();
 FILLCELL_X32 FILLCELL_70_384 ();
 FILLCELL_X32 FILLCELL_70_416 ();
 FILLCELL_X32 FILLCELL_70_448 ();
 FILLCELL_X32 FILLCELL_70_480 ();
 FILLCELL_X32 FILLCELL_70_512 ();
 FILLCELL_X32 FILLCELL_70_544 ();
 FILLCELL_X32 FILLCELL_70_576 ();
 FILLCELL_X32 FILLCELL_70_608 ();
 FILLCELL_X32 FILLCELL_70_640 ();
 FILLCELL_X32 FILLCELL_70_672 ();
 FILLCELL_X32 FILLCELL_70_704 ();
 FILLCELL_X32 FILLCELL_70_736 ();
 FILLCELL_X32 FILLCELL_70_768 ();
 FILLCELL_X32 FILLCELL_70_800 ();
 FILLCELL_X4 FILLCELL_70_832 ();
 FILLCELL_X32 FILLCELL_70_840 ();
 FILLCELL_X32 FILLCELL_70_872 ();
 FILLCELL_X32 FILLCELL_70_904 ();
 FILLCELL_X32 FILLCELL_70_936 ();
 FILLCELL_X32 FILLCELL_70_968 ();
 FILLCELL_X32 FILLCELL_70_1000 ();
 FILLCELL_X32 FILLCELL_70_1032 ();
 FILLCELL_X32 FILLCELL_70_1064 ();
 FILLCELL_X32 FILLCELL_70_1096 ();
 FILLCELL_X32 FILLCELL_70_1128 ();
 FILLCELL_X32 FILLCELL_70_1160 ();
 FILLCELL_X32 FILLCELL_70_1192 ();
 FILLCELL_X32 FILLCELL_70_1224 ();
 FILLCELL_X32 FILLCELL_70_1256 ();
 FILLCELL_X32 FILLCELL_70_1288 ();
 FILLCELL_X32 FILLCELL_70_1320 ();
 FILLCELL_X32 FILLCELL_70_1352 ();
 FILLCELL_X32 FILLCELL_70_1384 ();
 FILLCELL_X32 FILLCELL_70_1416 ();
 FILLCELL_X32 FILLCELL_70_1448 ();
 FILLCELL_X32 FILLCELL_70_1480 ();
 FILLCELL_X32 FILLCELL_70_1512 ();
 FILLCELL_X32 FILLCELL_70_1544 ();
 FILLCELL_X32 FILLCELL_70_1576 ();
 FILLCELL_X32 FILLCELL_70_1608 ();
 FILLCELL_X32 FILLCELL_70_1640 ();
 FILLCELL_X32 FILLCELL_70_1672 ();
 FILLCELL_X32 FILLCELL_70_1704 ();
 FILLCELL_X32 FILLCELL_70_1736 ();
 FILLCELL_X32 FILLCELL_70_1768 ();
 FILLCELL_X32 FILLCELL_70_1800 ();
 FILLCELL_X32 FILLCELL_70_1832 ();
 FILLCELL_X32 FILLCELL_70_1864 ();
 FILLCELL_X1 FILLCELL_70_1896 ();
 FILLCELL_X32 FILLCELL_71_0 ();
 FILLCELL_X32 FILLCELL_71_32 ();
 FILLCELL_X32 FILLCELL_71_64 ();
 FILLCELL_X32 FILLCELL_71_96 ();
 FILLCELL_X32 FILLCELL_71_128 ();
 FILLCELL_X32 FILLCELL_71_160 ();
 FILLCELL_X32 FILLCELL_71_192 ();
 FILLCELL_X32 FILLCELL_71_224 ();
 FILLCELL_X32 FILLCELL_71_256 ();
 FILLCELL_X32 FILLCELL_71_288 ();
 FILLCELL_X32 FILLCELL_71_320 ();
 FILLCELL_X32 FILLCELL_71_352 ();
 FILLCELL_X4 FILLCELL_71_384 ();
 FILLCELL_X2 FILLCELL_71_388 ();
 FILLCELL_X1 FILLCELL_71_390 ();
 FILLCELL_X32 FILLCELL_71_396 ();
 FILLCELL_X32 FILLCELL_71_428 ();
 FILLCELL_X16 FILLCELL_71_460 ();
 FILLCELL_X2 FILLCELL_71_476 ();
 FILLCELL_X1 FILLCELL_71_478 ();
 FILLCELL_X32 FILLCELL_71_484 ();
 FILLCELL_X32 FILLCELL_71_516 ();
 FILLCELL_X16 FILLCELL_71_548 ();
 FILLCELL_X32 FILLCELL_71_567 ();
 FILLCELL_X32 FILLCELL_71_599 ();
 FILLCELL_X32 FILLCELL_71_631 ();
 FILLCELL_X32 FILLCELL_71_663 ();
 FILLCELL_X16 FILLCELL_71_695 ();
 FILLCELL_X8 FILLCELL_71_711 ();
 FILLCELL_X16 FILLCELL_71_721 ();
 FILLCELL_X8 FILLCELL_71_737 ();
 FILLCELL_X2 FILLCELL_71_745 ();
 FILLCELL_X1 FILLCELL_71_747 ();
 FILLCELL_X32 FILLCELL_71_765 ();
 FILLCELL_X16 FILLCELL_71_797 ();
 FILLCELL_X8 FILLCELL_71_813 ();
 FILLCELL_X2 FILLCELL_71_821 ();
 FILLCELL_X1 FILLCELL_71_823 ();
 FILLCELL_X32 FILLCELL_71_829 ();
 FILLCELL_X32 FILLCELL_71_861 ();
 FILLCELL_X16 FILLCELL_71_893 ();
 FILLCELL_X32 FILLCELL_71_913 ();
 FILLCELL_X32 FILLCELL_71_945 ();
 FILLCELL_X32 FILLCELL_71_977 ();
 FILLCELL_X32 FILLCELL_71_1009 ();
 FILLCELL_X32 FILLCELL_71_1041 ();
 FILLCELL_X32 FILLCELL_71_1073 ();
 FILLCELL_X32 FILLCELL_71_1105 ();
 FILLCELL_X32 FILLCELL_71_1137 ();
 FILLCELL_X32 FILLCELL_71_1169 ();
 FILLCELL_X32 FILLCELL_71_1201 ();
 FILLCELL_X32 FILLCELL_71_1233 ();
 FILLCELL_X32 FILLCELL_71_1265 ();
 FILLCELL_X32 FILLCELL_71_1297 ();
 FILLCELL_X32 FILLCELL_71_1329 ();
 FILLCELL_X32 FILLCELL_71_1361 ();
 FILLCELL_X32 FILLCELL_71_1393 ();
 FILLCELL_X32 FILLCELL_71_1425 ();
 FILLCELL_X32 FILLCELL_71_1457 ();
 FILLCELL_X32 FILLCELL_71_1489 ();
 FILLCELL_X32 FILLCELL_71_1521 ();
 FILLCELL_X32 FILLCELL_71_1553 ();
 FILLCELL_X32 FILLCELL_71_1585 ();
 FILLCELL_X32 FILLCELL_71_1617 ();
 FILLCELL_X32 FILLCELL_71_1649 ();
 FILLCELL_X32 FILLCELL_71_1681 ();
 FILLCELL_X32 FILLCELL_71_1713 ();
 FILLCELL_X32 FILLCELL_71_1745 ();
 FILLCELL_X32 FILLCELL_71_1777 ();
 FILLCELL_X32 FILLCELL_71_1809 ();
 FILLCELL_X32 FILLCELL_71_1841 ();
 FILLCELL_X16 FILLCELL_71_1873 ();
 FILLCELL_X8 FILLCELL_71_1889 ();
 FILLCELL_X32 FILLCELL_72_0 ();
 FILLCELL_X32 FILLCELL_72_32 ();
 FILLCELL_X32 FILLCELL_72_64 ();
 FILLCELL_X32 FILLCELL_72_96 ();
 FILLCELL_X32 FILLCELL_72_128 ();
 FILLCELL_X32 FILLCELL_72_160 ();
 FILLCELL_X32 FILLCELL_72_192 ();
 FILLCELL_X32 FILLCELL_72_224 ();
 FILLCELL_X32 FILLCELL_72_256 ();
 FILLCELL_X32 FILLCELL_72_288 ();
 FILLCELL_X32 FILLCELL_72_320 ();
 FILLCELL_X32 FILLCELL_72_352 ();
 FILLCELL_X32 FILLCELL_72_384 ();
 FILLCELL_X32 FILLCELL_72_416 ();
 FILLCELL_X32 FILLCELL_72_448 ();
 FILLCELL_X32 FILLCELL_72_480 ();
 FILLCELL_X32 FILLCELL_72_512 ();
 FILLCELL_X32 FILLCELL_72_544 ();
 FILLCELL_X32 FILLCELL_72_576 ();
 FILLCELL_X32 FILLCELL_72_608 ();
 FILLCELL_X32 FILLCELL_72_640 ();
 FILLCELL_X32 FILLCELL_72_672 ();
 FILLCELL_X32 FILLCELL_72_704 ();
 FILLCELL_X32 FILLCELL_72_736 ();
 FILLCELL_X16 FILLCELL_72_768 ();
 FILLCELL_X4 FILLCELL_72_784 ();
 FILLCELL_X2 FILLCELL_72_788 ();
 FILLCELL_X32 FILLCELL_72_797 ();
 FILLCELL_X32 FILLCELL_72_829 ();
 FILLCELL_X32 FILLCELL_72_861 ();
 FILLCELL_X32 FILLCELL_72_893 ();
 FILLCELL_X1 FILLCELL_72_925 ();
 FILLCELL_X32 FILLCELL_72_930 ();
 FILLCELL_X32 FILLCELL_72_962 ();
 FILLCELL_X32 FILLCELL_72_994 ();
 FILLCELL_X32 FILLCELL_72_1026 ();
 FILLCELL_X32 FILLCELL_72_1058 ();
 FILLCELL_X32 FILLCELL_72_1090 ();
 FILLCELL_X32 FILLCELL_72_1122 ();
 FILLCELL_X32 FILLCELL_72_1154 ();
 FILLCELL_X32 FILLCELL_72_1186 ();
 FILLCELL_X32 FILLCELL_72_1218 ();
 FILLCELL_X32 FILLCELL_72_1250 ();
 FILLCELL_X32 FILLCELL_72_1282 ();
 FILLCELL_X32 FILLCELL_72_1314 ();
 FILLCELL_X32 FILLCELL_72_1346 ();
 FILLCELL_X32 FILLCELL_72_1378 ();
 FILLCELL_X32 FILLCELL_72_1410 ();
 FILLCELL_X32 FILLCELL_72_1442 ();
 FILLCELL_X32 FILLCELL_72_1474 ();
 FILLCELL_X32 FILLCELL_72_1506 ();
 FILLCELL_X32 FILLCELL_72_1538 ();
 FILLCELL_X32 FILLCELL_72_1570 ();
 FILLCELL_X32 FILLCELL_72_1602 ();
 FILLCELL_X32 FILLCELL_72_1634 ();
 FILLCELL_X32 FILLCELL_72_1666 ();
 FILLCELL_X32 FILLCELL_72_1698 ();
 FILLCELL_X32 FILLCELL_72_1730 ();
 FILLCELL_X32 FILLCELL_72_1762 ();
 FILLCELL_X32 FILLCELL_72_1794 ();
 FILLCELL_X32 FILLCELL_72_1826 ();
 FILLCELL_X32 FILLCELL_72_1858 ();
 FILLCELL_X4 FILLCELL_72_1890 ();
 FILLCELL_X2 FILLCELL_72_1894 ();
 FILLCELL_X1 FILLCELL_72_1896 ();
 FILLCELL_X32 FILLCELL_73_0 ();
 FILLCELL_X32 FILLCELL_73_32 ();
 FILLCELL_X32 FILLCELL_73_64 ();
 FILLCELL_X32 FILLCELL_73_96 ();
 FILLCELL_X32 FILLCELL_73_128 ();
 FILLCELL_X32 FILLCELL_73_160 ();
 FILLCELL_X32 FILLCELL_73_192 ();
 FILLCELL_X32 FILLCELL_73_224 ();
 FILLCELL_X32 FILLCELL_73_256 ();
 FILLCELL_X32 FILLCELL_73_288 ();
 FILLCELL_X32 FILLCELL_73_320 ();
 FILLCELL_X32 FILLCELL_73_352 ();
 FILLCELL_X32 FILLCELL_73_384 ();
 FILLCELL_X32 FILLCELL_73_416 ();
 FILLCELL_X32 FILLCELL_73_448 ();
 FILLCELL_X32 FILLCELL_73_480 ();
 FILLCELL_X32 FILLCELL_73_512 ();
 FILLCELL_X32 FILLCELL_73_544 ();
 FILLCELL_X32 FILLCELL_73_576 ();
 FILLCELL_X32 FILLCELL_73_608 ();
 FILLCELL_X32 FILLCELL_73_640 ();
 FILLCELL_X16 FILLCELL_73_672 ();
 FILLCELL_X8 FILLCELL_73_688 ();
 FILLCELL_X4 FILLCELL_73_696 ();
 FILLCELL_X1 FILLCELL_73_700 ();
 FILLCELL_X32 FILLCELL_73_704 ();
 FILLCELL_X32 FILLCELL_73_736 ();
 FILLCELL_X32 FILLCELL_73_768 ();
 FILLCELL_X32 FILLCELL_73_800 ();
 FILLCELL_X32 FILLCELL_73_832 ();
 FILLCELL_X32 FILLCELL_73_864 ();
 FILLCELL_X32 FILLCELL_73_896 ();
 FILLCELL_X4 FILLCELL_73_928 ();
 FILLCELL_X1 FILLCELL_73_932 ();
 FILLCELL_X32 FILLCELL_73_950 ();
 FILLCELL_X32 FILLCELL_73_982 ();
 FILLCELL_X32 FILLCELL_73_1014 ();
 FILLCELL_X32 FILLCELL_73_1046 ();
 FILLCELL_X32 FILLCELL_73_1078 ();
 FILLCELL_X32 FILLCELL_73_1110 ();
 FILLCELL_X32 FILLCELL_73_1142 ();
 FILLCELL_X32 FILLCELL_73_1174 ();
 FILLCELL_X32 FILLCELL_73_1206 ();
 FILLCELL_X32 FILLCELL_73_1238 ();
 FILLCELL_X32 FILLCELL_73_1270 ();
 FILLCELL_X32 FILLCELL_73_1302 ();
 FILLCELL_X32 FILLCELL_73_1334 ();
 FILLCELL_X32 FILLCELL_73_1366 ();
 FILLCELL_X32 FILLCELL_73_1398 ();
 FILLCELL_X32 FILLCELL_73_1430 ();
 FILLCELL_X32 FILLCELL_73_1462 ();
 FILLCELL_X32 FILLCELL_73_1494 ();
 FILLCELL_X32 FILLCELL_73_1526 ();
 FILLCELL_X32 FILLCELL_73_1558 ();
 FILLCELL_X32 FILLCELL_73_1590 ();
 FILLCELL_X32 FILLCELL_73_1622 ();
 FILLCELL_X32 FILLCELL_73_1654 ();
 FILLCELL_X32 FILLCELL_73_1686 ();
 FILLCELL_X32 FILLCELL_73_1718 ();
 FILLCELL_X32 FILLCELL_73_1750 ();
 FILLCELL_X32 FILLCELL_73_1782 ();
 FILLCELL_X32 FILLCELL_73_1814 ();
 FILLCELL_X32 FILLCELL_73_1846 ();
 FILLCELL_X16 FILLCELL_73_1878 ();
 FILLCELL_X2 FILLCELL_73_1894 ();
 FILLCELL_X1 FILLCELL_73_1896 ();
 FILLCELL_X32 FILLCELL_74_0 ();
 FILLCELL_X32 FILLCELL_74_32 ();
 FILLCELL_X32 FILLCELL_74_64 ();
 FILLCELL_X32 FILLCELL_74_96 ();
 FILLCELL_X4 FILLCELL_74_128 ();
 FILLCELL_X32 FILLCELL_74_149 ();
 FILLCELL_X32 FILLCELL_74_181 ();
 FILLCELL_X32 FILLCELL_74_213 ();
 FILLCELL_X32 FILLCELL_74_245 ();
 FILLCELL_X16 FILLCELL_74_277 ();
 FILLCELL_X4 FILLCELL_74_293 ();
 FILLCELL_X2 FILLCELL_74_297 ();
 FILLCELL_X1 FILLCELL_74_299 ();
 FILLCELL_X32 FILLCELL_74_302 ();
 FILLCELL_X32 FILLCELL_74_334 ();
 FILLCELL_X32 FILLCELL_74_366 ();
 FILLCELL_X16 FILLCELL_74_398 ();
 FILLCELL_X2 FILLCELL_74_414 ();
 FILLCELL_X32 FILLCELL_74_419 ();
 FILLCELL_X32 FILLCELL_74_451 ();
 FILLCELL_X32 FILLCELL_74_483 ();
 FILLCELL_X32 FILLCELL_74_515 ();
 FILLCELL_X32 FILLCELL_74_547 ();
 FILLCELL_X8 FILLCELL_74_579 ();
 FILLCELL_X4 FILLCELL_74_587 ();
 FILLCELL_X2 FILLCELL_74_591 ();
 FILLCELL_X32 FILLCELL_74_598 ();
 FILLCELL_X32 FILLCELL_74_630 ();
 FILLCELL_X32 FILLCELL_74_662 ();
 FILLCELL_X8 FILLCELL_74_694 ();
 FILLCELL_X32 FILLCELL_74_705 ();
 FILLCELL_X32 FILLCELL_74_737 ();
 FILLCELL_X32 FILLCELL_74_769 ();
 FILLCELL_X32 FILLCELL_74_801 ();
 FILLCELL_X8 FILLCELL_74_833 ();
 FILLCELL_X2 FILLCELL_74_841 ();
 FILLCELL_X32 FILLCELL_74_846 ();
 FILLCELL_X32 FILLCELL_74_878 ();
 FILLCELL_X16 FILLCELL_74_910 ();
 FILLCELL_X2 FILLCELL_74_926 ();
 FILLCELL_X32 FILLCELL_74_931 ();
 FILLCELL_X32 FILLCELL_74_963 ();
 FILLCELL_X32 FILLCELL_74_995 ();
 FILLCELL_X32 FILLCELL_74_1027 ();
 FILLCELL_X32 FILLCELL_74_1059 ();
 FILLCELL_X32 FILLCELL_74_1091 ();
 FILLCELL_X32 FILLCELL_74_1123 ();
 FILLCELL_X32 FILLCELL_74_1155 ();
 FILLCELL_X32 FILLCELL_74_1187 ();
 FILLCELL_X32 FILLCELL_74_1219 ();
 FILLCELL_X32 FILLCELL_74_1251 ();
 FILLCELL_X32 FILLCELL_74_1283 ();
 FILLCELL_X32 FILLCELL_74_1315 ();
 FILLCELL_X32 FILLCELL_74_1347 ();
 FILLCELL_X32 FILLCELL_74_1379 ();
 FILLCELL_X32 FILLCELL_74_1411 ();
 FILLCELL_X32 FILLCELL_74_1443 ();
 FILLCELL_X32 FILLCELL_74_1475 ();
 FILLCELL_X32 FILLCELL_74_1507 ();
 FILLCELL_X32 FILLCELL_74_1539 ();
 FILLCELL_X32 FILLCELL_74_1571 ();
 FILLCELL_X32 FILLCELL_74_1603 ();
 FILLCELL_X32 FILLCELL_74_1635 ();
 FILLCELL_X32 FILLCELL_74_1667 ();
 FILLCELL_X32 FILLCELL_74_1699 ();
 FILLCELL_X32 FILLCELL_74_1731 ();
 FILLCELL_X32 FILLCELL_74_1763 ();
 FILLCELL_X32 FILLCELL_74_1795 ();
 FILLCELL_X32 FILLCELL_74_1827 ();
 FILLCELL_X32 FILLCELL_74_1859 ();
 FILLCELL_X4 FILLCELL_74_1891 ();
 FILLCELL_X2 FILLCELL_74_1895 ();
 FILLCELL_X32 FILLCELL_75_0 ();
 FILLCELL_X32 FILLCELL_75_32 ();
 FILLCELL_X32 FILLCELL_75_64 ();
 FILLCELL_X32 FILLCELL_75_96 ();
 FILLCELL_X32 FILLCELL_75_128 ();
 FILLCELL_X32 FILLCELL_75_160 ();
 FILLCELL_X32 FILLCELL_75_192 ();
 FILLCELL_X32 FILLCELL_75_224 ();
 FILLCELL_X32 FILLCELL_75_256 ();
 FILLCELL_X32 FILLCELL_75_288 ();
 FILLCELL_X32 FILLCELL_75_320 ();
 FILLCELL_X32 FILLCELL_75_352 ();
 FILLCELL_X32 FILLCELL_75_384 ();
 FILLCELL_X32 FILLCELL_75_416 ();
 FILLCELL_X32 FILLCELL_75_448 ();
 FILLCELL_X32 FILLCELL_75_480 ();
 FILLCELL_X32 FILLCELL_75_512 ();
 FILLCELL_X32 FILLCELL_75_544 ();
 FILLCELL_X16 FILLCELL_75_576 ();
 FILLCELL_X32 FILLCELL_75_595 ();
 FILLCELL_X32 FILLCELL_75_627 ();
 FILLCELL_X16 FILLCELL_75_659 ();
 FILLCELL_X8 FILLCELL_75_675 ();
 FILLCELL_X4 FILLCELL_75_683 ();
 FILLCELL_X32 FILLCELL_75_691 ();
 FILLCELL_X8 FILLCELL_75_723 ();
 FILLCELL_X4 FILLCELL_75_731 ();
 FILLCELL_X2 FILLCELL_75_735 ();
 FILLCELL_X1 FILLCELL_75_737 ();
 FILLCELL_X32 FILLCELL_75_740 ();
 FILLCELL_X32 FILLCELL_75_772 ();
 FILLCELL_X32 FILLCELL_75_804 ();
 FILLCELL_X32 FILLCELL_75_836 ();
 FILLCELL_X32 FILLCELL_75_868 ();
 FILLCELL_X32 FILLCELL_75_900 ();
 FILLCELL_X32 FILLCELL_75_932 ();
 FILLCELL_X32 FILLCELL_75_964 ();
 FILLCELL_X32 FILLCELL_75_996 ();
 FILLCELL_X32 FILLCELL_75_1028 ();
 FILLCELL_X32 FILLCELL_75_1060 ();
 FILLCELL_X32 FILLCELL_75_1092 ();
 FILLCELL_X32 FILLCELL_75_1124 ();
 FILLCELL_X32 FILLCELL_75_1156 ();
 FILLCELL_X32 FILLCELL_75_1188 ();
 FILLCELL_X32 FILLCELL_75_1220 ();
 FILLCELL_X32 FILLCELL_75_1252 ();
 FILLCELL_X32 FILLCELL_75_1284 ();
 FILLCELL_X32 FILLCELL_75_1316 ();
 FILLCELL_X32 FILLCELL_75_1348 ();
 FILLCELL_X32 FILLCELL_75_1380 ();
 FILLCELL_X32 FILLCELL_75_1412 ();
 FILLCELL_X32 FILLCELL_75_1444 ();
 FILLCELL_X32 FILLCELL_75_1476 ();
 FILLCELL_X32 FILLCELL_75_1508 ();
 FILLCELL_X32 FILLCELL_75_1540 ();
 FILLCELL_X32 FILLCELL_75_1572 ();
 FILLCELL_X32 FILLCELL_75_1604 ();
 FILLCELL_X32 FILLCELL_75_1636 ();
 FILLCELL_X32 FILLCELL_75_1668 ();
 FILLCELL_X32 FILLCELL_75_1700 ();
 FILLCELL_X32 FILLCELL_75_1732 ();
 FILLCELL_X32 FILLCELL_75_1764 ();
 FILLCELL_X32 FILLCELL_75_1796 ();
 FILLCELL_X32 FILLCELL_75_1828 ();
 FILLCELL_X32 FILLCELL_75_1860 ();
 FILLCELL_X4 FILLCELL_75_1892 ();
 FILLCELL_X1 FILLCELL_75_1896 ();
 FILLCELL_X32 FILLCELL_76_0 ();
 FILLCELL_X32 FILLCELL_76_32 ();
 FILLCELL_X32 FILLCELL_76_64 ();
 FILLCELL_X32 FILLCELL_76_96 ();
 FILLCELL_X32 FILLCELL_76_128 ();
 FILLCELL_X32 FILLCELL_76_160 ();
 FILLCELL_X16 FILLCELL_76_192 ();
 FILLCELL_X32 FILLCELL_76_212 ();
 FILLCELL_X32 FILLCELL_76_244 ();
 FILLCELL_X16 FILLCELL_76_276 ();
 FILLCELL_X8 FILLCELL_76_292 ();
 FILLCELL_X1 FILLCELL_76_300 ();
 FILLCELL_X4 FILLCELL_76_304 ();
 FILLCELL_X2 FILLCELL_76_308 ();
 FILLCELL_X1 FILLCELL_76_310 ();
 FILLCELL_X32 FILLCELL_76_316 ();
 FILLCELL_X32 FILLCELL_76_348 ();
 FILLCELL_X16 FILLCELL_76_380 ();
 FILLCELL_X32 FILLCELL_76_400 ();
 FILLCELL_X32 FILLCELL_76_432 ();
 FILLCELL_X32 FILLCELL_76_464 ();
 FILLCELL_X32 FILLCELL_76_496 ();
 FILLCELL_X32 FILLCELL_76_528 ();
 FILLCELL_X32 FILLCELL_76_560 ();
 FILLCELL_X32 FILLCELL_76_592 ();
 FILLCELL_X32 FILLCELL_76_624 ();
 FILLCELL_X2 FILLCELL_76_656 ();
 FILLCELL_X32 FILLCELL_76_661 ();
 FILLCELL_X32 FILLCELL_76_693 ();
 FILLCELL_X32 FILLCELL_76_725 ();
 FILLCELL_X32 FILLCELL_76_757 ();
 FILLCELL_X32 FILLCELL_76_789 ();
 FILLCELL_X32 FILLCELL_76_821 ();
 FILLCELL_X32 FILLCELL_76_853 ();
 FILLCELL_X32 FILLCELL_76_885 ();
 FILLCELL_X32 FILLCELL_76_917 ();
 FILLCELL_X32 FILLCELL_76_949 ();
 FILLCELL_X32 FILLCELL_76_981 ();
 FILLCELL_X16 FILLCELL_76_1013 ();
 FILLCELL_X8 FILLCELL_76_1029 ();
 FILLCELL_X4 FILLCELL_76_1037 ();
 FILLCELL_X32 FILLCELL_76_1043 ();
 FILLCELL_X32 FILLCELL_76_1075 ();
 FILLCELL_X32 FILLCELL_76_1107 ();
 FILLCELL_X32 FILLCELL_76_1139 ();
 FILLCELL_X32 FILLCELL_76_1171 ();
 FILLCELL_X32 FILLCELL_76_1203 ();
 FILLCELL_X32 FILLCELL_76_1235 ();
 FILLCELL_X32 FILLCELL_76_1267 ();
 FILLCELL_X32 FILLCELL_76_1299 ();
 FILLCELL_X32 FILLCELL_76_1331 ();
 FILLCELL_X32 FILLCELL_76_1363 ();
 FILLCELL_X32 FILLCELL_76_1395 ();
 FILLCELL_X32 FILLCELL_76_1427 ();
 FILLCELL_X32 FILLCELL_76_1459 ();
 FILLCELL_X32 FILLCELL_76_1491 ();
 FILLCELL_X32 FILLCELL_76_1523 ();
 FILLCELL_X32 FILLCELL_76_1555 ();
 FILLCELL_X32 FILLCELL_76_1587 ();
 FILLCELL_X32 FILLCELL_76_1619 ();
 FILLCELL_X32 FILLCELL_76_1651 ();
 FILLCELL_X32 FILLCELL_76_1683 ();
 FILLCELL_X32 FILLCELL_76_1715 ();
 FILLCELL_X32 FILLCELL_76_1747 ();
 FILLCELL_X32 FILLCELL_76_1779 ();
 FILLCELL_X32 FILLCELL_76_1811 ();
 FILLCELL_X32 FILLCELL_76_1843 ();
 FILLCELL_X16 FILLCELL_76_1875 ();
 FILLCELL_X4 FILLCELL_76_1891 ();
 FILLCELL_X2 FILLCELL_76_1895 ();
 FILLCELL_X32 FILLCELL_77_0 ();
 FILLCELL_X32 FILLCELL_77_32 ();
 FILLCELL_X32 FILLCELL_77_64 ();
 FILLCELL_X32 FILLCELL_77_96 ();
 FILLCELL_X32 FILLCELL_77_128 ();
 FILLCELL_X32 FILLCELL_77_160 ();
 FILLCELL_X8 FILLCELL_77_192 ();
 FILLCELL_X4 FILLCELL_77_200 ();
 FILLCELL_X1 FILLCELL_77_204 ();
 FILLCELL_X32 FILLCELL_77_208 ();
 FILLCELL_X32 FILLCELL_77_240 ();
 FILLCELL_X32 FILLCELL_77_272 ();
 FILLCELL_X32 FILLCELL_77_304 ();
 FILLCELL_X32 FILLCELL_77_336 ();
 FILLCELL_X16 FILLCELL_77_368 ();
 FILLCELL_X8 FILLCELL_77_384 ();
 FILLCELL_X4 FILLCELL_77_392 ();
 FILLCELL_X2 FILLCELL_77_396 ();
 FILLCELL_X32 FILLCELL_77_401 ();
 FILLCELL_X32 FILLCELL_77_433 ();
 FILLCELL_X32 FILLCELL_77_465 ();
 FILLCELL_X32 FILLCELL_77_497 ();
 FILLCELL_X32 FILLCELL_77_529 ();
 FILLCELL_X32 FILLCELL_77_561 ();
 FILLCELL_X16 FILLCELL_77_593 ();
 FILLCELL_X8 FILLCELL_77_609 ();
 FILLCELL_X4 FILLCELL_77_617 ();
 FILLCELL_X32 FILLCELL_77_625 ();
 FILLCELL_X32 FILLCELL_77_657 ();
 FILLCELL_X32 FILLCELL_77_689 ();
 FILLCELL_X32 FILLCELL_77_721 ();
 FILLCELL_X32 FILLCELL_77_753 ();
 FILLCELL_X32 FILLCELL_77_785 ();
 FILLCELL_X32 FILLCELL_77_817 ();
 FILLCELL_X32 FILLCELL_77_849 ();
 FILLCELL_X32 FILLCELL_77_881 ();
 FILLCELL_X32 FILLCELL_77_913 ();
 FILLCELL_X32 FILLCELL_77_945 ();
 FILLCELL_X32 FILLCELL_77_977 ();
 FILLCELL_X32 FILLCELL_77_1009 ();
 FILLCELL_X32 FILLCELL_77_1041 ();
 FILLCELL_X32 FILLCELL_77_1073 ();
 FILLCELL_X32 FILLCELL_77_1105 ();
 FILLCELL_X32 FILLCELL_77_1137 ();
 FILLCELL_X32 FILLCELL_77_1169 ();
 FILLCELL_X32 FILLCELL_77_1201 ();
 FILLCELL_X32 FILLCELL_77_1233 ();
 FILLCELL_X32 FILLCELL_77_1265 ();
 FILLCELL_X32 FILLCELL_77_1297 ();
 FILLCELL_X32 FILLCELL_77_1329 ();
 FILLCELL_X32 FILLCELL_77_1361 ();
 FILLCELL_X32 FILLCELL_77_1393 ();
 FILLCELL_X32 FILLCELL_77_1425 ();
 FILLCELL_X32 FILLCELL_77_1457 ();
 FILLCELL_X32 FILLCELL_77_1489 ();
 FILLCELL_X32 FILLCELL_77_1521 ();
 FILLCELL_X32 FILLCELL_77_1553 ();
 FILLCELL_X32 FILLCELL_77_1585 ();
 FILLCELL_X32 FILLCELL_77_1617 ();
 FILLCELL_X32 FILLCELL_77_1649 ();
 FILLCELL_X32 FILLCELL_77_1681 ();
 FILLCELL_X32 FILLCELL_77_1713 ();
 FILLCELL_X32 FILLCELL_77_1745 ();
 FILLCELL_X32 FILLCELL_77_1777 ();
 FILLCELL_X32 FILLCELL_77_1809 ();
 FILLCELL_X32 FILLCELL_77_1841 ();
 FILLCELL_X16 FILLCELL_77_1873 ();
 FILLCELL_X8 FILLCELL_77_1889 ();
 FILLCELL_X32 FILLCELL_78_0 ();
 FILLCELL_X32 FILLCELL_78_32 ();
 FILLCELL_X32 FILLCELL_78_64 ();
 FILLCELL_X32 FILLCELL_78_96 ();
 FILLCELL_X32 FILLCELL_78_128 ();
 FILLCELL_X32 FILLCELL_78_160 ();
 FILLCELL_X16 FILLCELL_78_192 ();
 FILLCELL_X8 FILLCELL_78_208 ();
 FILLCELL_X1 FILLCELL_78_216 ();
 FILLCELL_X4 FILLCELL_78_221 ();
 FILLCELL_X1 FILLCELL_78_225 ();
 FILLCELL_X16 FILLCELL_78_229 ();
 FILLCELL_X8 FILLCELL_78_245 ();
 FILLCELL_X2 FILLCELL_78_253 ();
 FILLCELL_X32 FILLCELL_78_259 ();
 FILLCELL_X32 FILLCELL_78_291 ();
 FILLCELL_X32 FILLCELL_78_323 ();
 FILLCELL_X32 FILLCELL_78_355 ();
 FILLCELL_X32 FILLCELL_78_387 ();
 FILLCELL_X32 FILLCELL_78_419 ();
 FILLCELL_X32 FILLCELL_78_451 ();
 FILLCELL_X32 FILLCELL_78_483 ();
 FILLCELL_X32 FILLCELL_78_515 ();
 FILLCELL_X32 FILLCELL_78_547 ();
 FILLCELL_X32 FILLCELL_78_579 ();
 FILLCELL_X32 FILLCELL_78_611 ();
 FILLCELL_X32 FILLCELL_78_643 ();
 FILLCELL_X32 FILLCELL_78_675 ();
 FILLCELL_X32 FILLCELL_78_707 ();
 FILLCELL_X32 FILLCELL_78_739 ();
 FILLCELL_X32 FILLCELL_78_771 ();
 FILLCELL_X32 FILLCELL_78_803 ();
 FILLCELL_X32 FILLCELL_78_835 ();
 FILLCELL_X32 FILLCELL_78_867 ();
 FILLCELL_X32 FILLCELL_78_899 ();
 FILLCELL_X32 FILLCELL_78_931 ();
 FILLCELL_X32 FILLCELL_78_963 ();
 FILLCELL_X32 FILLCELL_78_995 ();
 FILLCELL_X32 FILLCELL_78_1027 ();
 FILLCELL_X32 FILLCELL_78_1059 ();
 FILLCELL_X32 FILLCELL_78_1091 ();
 FILLCELL_X32 FILLCELL_78_1123 ();
 FILLCELL_X32 FILLCELL_78_1155 ();
 FILLCELL_X32 FILLCELL_78_1187 ();
 FILLCELL_X32 FILLCELL_78_1219 ();
 FILLCELL_X32 FILLCELL_78_1251 ();
 FILLCELL_X32 FILLCELL_78_1283 ();
 FILLCELL_X32 FILLCELL_78_1315 ();
 FILLCELL_X32 FILLCELL_78_1347 ();
 FILLCELL_X32 FILLCELL_78_1379 ();
 FILLCELL_X32 FILLCELL_78_1411 ();
 FILLCELL_X32 FILLCELL_78_1443 ();
 FILLCELL_X32 FILLCELL_78_1475 ();
 FILLCELL_X32 FILLCELL_78_1507 ();
 FILLCELL_X32 FILLCELL_78_1539 ();
 FILLCELL_X32 FILLCELL_78_1571 ();
 FILLCELL_X32 FILLCELL_78_1603 ();
 FILLCELL_X32 FILLCELL_78_1635 ();
 FILLCELL_X32 FILLCELL_78_1667 ();
 FILLCELL_X32 FILLCELL_78_1699 ();
 FILLCELL_X32 FILLCELL_78_1731 ();
 FILLCELL_X32 FILLCELL_78_1763 ();
 FILLCELL_X32 FILLCELL_78_1795 ();
 FILLCELL_X32 FILLCELL_78_1827 ();
 FILLCELL_X32 FILLCELL_78_1859 ();
 FILLCELL_X4 FILLCELL_78_1891 ();
 FILLCELL_X2 FILLCELL_78_1895 ();
 FILLCELL_X32 FILLCELL_79_0 ();
 FILLCELL_X32 FILLCELL_79_32 ();
 FILLCELL_X32 FILLCELL_79_64 ();
 FILLCELL_X32 FILLCELL_79_96 ();
 FILLCELL_X32 FILLCELL_79_128 ();
 FILLCELL_X32 FILLCELL_79_160 ();
 FILLCELL_X32 FILLCELL_79_192 ();
 FILLCELL_X16 FILLCELL_79_224 ();
 FILLCELL_X4 FILLCELL_79_240 ();
 FILLCELL_X32 FILLCELL_79_247 ();
 FILLCELL_X32 FILLCELL_79_279 ();
 FILLCELL_X32 FILLCELL_79_311 ();
 FILLCELL_X32 FILLCELL_79_343 ();
 FILLCELL_X32 FILLCELL_79_375 ();
 FILLCELL_X32 FILLCELL_79_407 ();
 FILLCELL_X32 FILLCELL_79_439 ();
 FILLCELL_X32 FILLCELL_79_471 ();
 FILLCELL_X32 FILLCELL_79_503 ();
 FILLCELL_X4 FILLCELL_79_535 ();
 FILLCELL_X32 FILLCELL_79_543 ();
 FILLCELL_X32 FILLCELL_79_575 ();
 FILLCELL_X32 FILLCELL_79_607 ();
 FILLCELL_X32 FILLCELL_79_639 ();
 FILLCELL_X32 FILLCELL_79_671 ();
 FILLCELL_X32 FILLCELL_79_703 ();
 FILLCELL_X32 FILLCELL_79_735 ();
 FILLCELL_X32 FILLCELL_79_767 ();
 FILLCELL_X32 FILLCELL_79_799 ();
 FILLCELL_X32 FILLCELL_79_831 ();
 FILLCELL_X32 FILLCELL_79_863 ();
 FILLCELL_X32 FILLCELL_79_895 ();
 FILLCELL_X32 FILLCELL_79_927 ();
 FILLCELL_X32 FILLCELL_79_959 ();
 FILLCELL_X32 FILLCELL_79_991 ();
 FILLCELL_X16 FILLCELL_79_1023 ();
 FILLCELL_X8 FILLCELL_79_1039 ();
 FILLCELL_X4 FILLCELL_79_1047 ();
 FILLCELL_X2 FILLCELL_79_1051 ();
 FILLCELL_X32 FILLCELL_79_1070 ();
 FILLCELL_X32 FILLCELL_79_1102 ();
 FILLCELL_X32 FILLCELL_79_1134 ();
 FILLCELL_X32 FILLCELL_79_1166 ();
 FILLCELL_X32 FILLCELL_79_1198 ();
 FILLCELL_X32 FILLCELL_79_1230 ();
 FILLCELL_X32 FILLCELL_79_1262 ();
 FILLCELL_X32 FILLCELL_79_1294 ();
 FILLCELL_X32 FILLCELL_79_1326 ();
 FILLCELL_X32 FILLCELL_79_1358 ();
 FILLCELL_X32 FILLCELL_79_1390 ();
 FILLCELL_X32 FILLCELL_79_1422 ();
 FILLCELL_X32 FILLCELL_79_1454 ();
 FILLCELL_X32 FILLCELL_79_1486 ();
 FILLCELL_X32 FILLCELL_79_1518 ();
 FILLCELL_X32 FILLCELL_79_1550 ();
 FILLCELL_X32 FILLCELL_79_1582 ();
 FILLCELL_X32 FILLCELL_79_1614 ();
 FILLCELL_X32 FILLCELL_79_1646 ();
 FILLCELL_X32 FILLCELL_79_1678 ();
 FILLCELL_X32 FILLCELL_79_1710 ();
 FILLCELL_X32 FILLCELL_79_1742 ();
 FILLCELL_X32 FILLCELL_79_1774 ();
 FILLCELL_X32 FILLCELL_79_1806 ();
 FILLCELL_X32 FILLCELL_79_1838 ();
 FILLCELL_X16 FILLCELL_79_1870 ();
 FILLCELL_X8 FILLCELL_79_1886 ();
 FILLCELL_X2 FILLCELL_79_1894 ();
 FILLCELL_X1 FILLCELL_79_1896 ();
 FILLCELL_X32 FILLCELL_80_0 ();
 FILLCELL_X32 FILLCELL_80_32 ();
 FILLCELL_X32 FILLCELL_80_64 ();
 FILLCELL_X32 FILLCELL_80_96 ();
 FILLCELL_X32 FILLCELL_80_128 ();
 FILLCELL_X32 FILLCELL_80_160 ();
 FILLCELL_X32 FILLCELL_80_192 ();
 FILLCELL_X32 FILLCELL_80_224 ();
 FILLCELL_X32 FILLCELL_80_256 ();
 FILLCELL_X16 FILLCELL_80_288 ();
 FILLCELL_X8 FILLCELL_80_304 ();
 FILLCELL_X4 FILLCELL_80_312 ();
 FILLCELL_X32 FILLCELL_80_321 ();
 FILLCELL_X32 FILLCELL_80_353 ();
 FILLCELL_X1 FILLCELL_80_385 ();
 FILLCELL_X32 FILLCELL_80_389 ();
 FILLCELL_X32 FILLCELL_80_421 ();
 FILLCELL_X32 FILLCELL_80_453 ();
 FILLCELL_X32 FILLCELL_80_485 ();
 FILLCELL_X32 FILLCELL_80_517 ();
 FILLCELL_X4 FILLCELL_80_549 ();
 FILLCELL_X32 FILLCELL_80_555 ();
 FILLCELL_X32 FILLCELL_80_587 ();
 FILLCELL_X32 FILLCELL_80_619 ();
 FILLCELL_X32 FILLCELL_80_651 ();
 FILLCELL_X32 FILLCELL_80_683 ();
 FILLCELL_X32 FILLCELL_80_715 ();
 FILLCELL_X32 FILLCELL_80_747 ();
 FILLCELL_X32 FILLCELL_80_779 ();
 FILLCELL_X32 FILLCELL_80_811 ();
 FILLCELL_X32 FILLCELL_80_843 ();
 FILLCELL_X32 FILLCELL_80_875 ();
 FILLCELL_X32 FILLCELL_80_907 ();
 FILLCELL_X32 FILLCELL_80_939 ();
 FILLCELL_X32 FILLCELL_80_971 ();
 FILLCELL_X32 FILLCELL_80_1003 ();
 FILLCELL_X1 FILLCELL_80_1035 ();
 FILLCELL_X32 FILLCELL_80_1043 ();
 FILLCELL_X32 FILLCELL_80_1075 ();
 FILLCELL_X32 FILLCELL_80_1107 ();
 FILLCELL_X32 FILLCELL_80_1139 ();
 FILLCELL_X32 FILLCELL_80_1171 ();
 FILLCELL_X32 FILLCELL_80_1203 ();
 FILLCELL_X32 FILLCELL_80_1235 ();
 FILLCELL_X32 FILLCELL_80_1267 ();
 FILLCELL_X32 FILLCELL_80_1299 ();
 FILLCELL_X32 FILLCELL_80_1331 ();
 FILLCELL_X32 FILLCELL_80_1363 ();
 FILLCELL_X32 FILLCELL_80_1395 ();
 FILLCELL_X32 FILLCELL_80_1427 ();
 FILLCELL_X32 FILLCELL_80_1459 ();
 FILLCELL_X32 FILLCELL_80_1491 ();
 FILLCELL_X32 FILLCELL_80_1523 ();
 FILLCELL_X32 FILLCELL_80_1555 ();
 FILLCELL_X32 FILLCELL_80_1587 ();
 FILLCELL_X32 FILLCELL_80_1619 ();
 FILLCELL_X32 FILLCELL_80_1651 ();
 FILLCELL_X32 FILLCELL_80_1683 ();
 FILLCELL_X32 FILLCELL_80_1715 ();
 FILLCELL_X32 FILLCELL_80_1747 ();
 FILLCELL_X32 FILLCELL_80_1779 ();
 FILLCELL_X32 FILLCELL_80_1811 ();
 FILLCELL_X32 FILLCELL_80_1843 ();
 FILLCELL_X16 FILLCELL_80_1875 ();
 FILLCELL_X4 FILLCELL_80_1891 ();
 FILLCELL_X2 FILLCELL_80_1895 ();
 FILLCELL_X32 FILLCELL_81_0 ();
 FILLCELL_X32 FILLCELL_81_32 ();
 FILLCELL_X32 FILLCELL_81_64 ();
 FILLCELL_X32 FILLCELL_81_96 ();
 FILLCELL_X32 FILLCELL_81_128 ();
 FILLCELL_X32 FILLCELL_81_160 ();
 FILLCELL_X32 FILLCELL_81_192 ();
 FILLCELL_X32 FILLCELL_81_224 ();
 FILLCELL_X32 FILLCELL_81_256 ();
 FILLCELL_X32 FILLCELL_81_288 ();
 FILLCELL_X32 FILLCELL_81_320 ();
 FILLCELL_X32 FILLCELL_81_352 ();
 FILLCELL_X32 FILLCELL_81_384 ();
 FILLCELL_X32 FILLCELL_81_416 ();
 FILLCELL_X32 FILLCELL_81_448 ();
 FILLCELL_X32 FILLCELL_81_480 ();
 FILLCELL_X32 FILLCELL_81_512 ();
 FILLCELL_X32 FILLCELL_81_544 ();
 FILLCELL_X32 FILLCELL_81_576 ();
 FILLCELL_X16 FILLCELL_81_608 ();
 FILLCELL_X4 FILLCELL_81_624 ();
 FILLCELL_X1 FILLCELL_81_628 ();
 FILLCELL_X32 FILLCELL_81_632 ();
 FILLCELL_X32 FILLCELL_81_664 ();
 FILLCELL_X32 FILLCELL_81_696 ();
 FILLCELL_X32 FILLCELL_81_728 ();
 FILLCELL_X32 FILLCELL_81_760 ();
 FILLCELL_X32 FILLCELL_81_792 ();
 FILLCELL_X32 FILLCELL_81_824 ();
 FILLCELL_X32 FILLCELL_81_856 ();
 FILLCELL_X32 FILLCELL_81_888 ();
 FILLCELL_X32 FILLCELL_81_920 ();
 FILLCELL_X32 FILLCELL_81_952 ();
 FILLCELL_X32 FILLCELL_81_984 ();
 FILLCELL_X16 FILLCELL_81_1016 ();
 FILLCELL_X4 FILLCELL_81_1032 ();
 FILLCELL_X2 FILLCELL_81_1036 ();
 FILLCELL_X32 FILLCELL_81_1042 ();
 FILLCELL_X32 FILLCELL_81_1074 ();
 FILLCELL_X32 FILLCELL_81_1106 ();
 FILLCELL_X32 FILLCELL_81_1138 ();
 FILLCELL_X32 FILLCELL_81_1170 ();
 FILLCELL_X32 FILLCELL_81_1202 ();
 FILLCELL_X32 FILLCELL_81_1234 ();
 FILLCELL_X32 FILLCELL_81_1266 ();
 FILLCELL_X32 FILLCELL_81_1298 ();
 FILLCELL_X32 FILLCELL_81_1330 ();
 FILLCELL_X32 FILLCELL_81_1362 ();
 FILLCELL_X32 FILLCELL_81_1394 ();
 FILLCELL_X32 FILLCELL_81_1426 ();
 FILLCELL_X32 FILLCELL_81_1458 ();
 FILLCELL_X32 FILLCELL_81_1490 ();
 FILLCELL_X32 FILLCELL_81_1522 ();
 FILLCELL_X32 FILLCELL_81_1554 ();
 FILLCELL_X32 FILLCELL_81_1586 ();
 FILLCELL_X32 FILLCELL_81_1618 ();
 FILLCELL_X32 FILLCELL_81_1650 ();
 FILLCELL_X32 FILLCELL_81_1682 ();
 FILLCELL_X32 FILLCELL_81_1714 ();
 FILLCELL_X32 FILLCELL_81_1746 ();
 FILLCELL_X32 FILLCELL_81_1778 ();
 FILLCELL_X32 FILLCELL_81_1810 ();
 FILLCELL_X32 FILLCELL_81_1842 ();
 FILLCELL_X16 FILLCELL_81_1874 ();
 FILLCELL_X4 FILLCELL_81_1890 ();
 FILLCELL_X2 FILLCELL_81_1894 ();
 FILLCELL_X1 FILLCELL_81_1896 ();
 FILLCELL_X32 FILLCELL_82_0 ();
 FILLCELL_X32 FILLCELL_82_32 ();
 FILLCELL_X32 FILLCELL_82_64 ();
 FILLCELL_X32 FILLCELL_82_96 ();
 FILLCELL_X32 FILLCELL_82_128 ();
 FILLCELL_X32 FILLCELL_82_160 ();
 FILLCELL_X32 FILLCELL_82_192 ();
 FILLCELL_X32 FILLCELL_82_224 ();
 FILLCELL_X32 FILLCELL_82_256 ();
 FILLCELL_X32 FILLCELL_82_288 ();
 FILLCELL_X32 FILLCELL_82_320 ();
 FILLCELL_X32 FILLCELL_82_352 ();
 FILLCELL_X32 FILLCELL_82_384 ();
 FILLCELL_X32 FILLCELL_82_416 ();
 FILLCELL_X8 FILLCELL_82_448 ();
 FILLCELL_X2 FILLCELL_82_456 ();
 FILLCELL_X16 FILLCELL_82_467 ();
 FILLCELL_X4 FILLCELL_82_483 ();
 FILLCELL_X2 FILLCELL_82_487 ();
 FILLCELL_X32 FILLCELL_82_491 ();
 FILLCELL_X32 FILLCELL_82_523 ();
 FILLCELL_X32 FILLCELL_82_560 ();
 FILLCELL_X32 FILLCELL_82_592 ();
 FILLCELL_X32 FILLCELL_82_624 ();
 FILLCELL_X16 FILLCELL_82_656 ();
 FILLCELL_X4 FILLCELL_82_672 ();
 FILLCELL_X1 FILLCELL_82_676 ();
 FILLCELL_X32 FILLCELL_82_680 ();
 FILLCELL_X32 FILLCELL_82_712 ();
 FILLCELL_X32 FILLCELL_82_744 ();
 FILLCELL_X32 FILLCELL_82_776 ();
 FILLCELL_X32 FILLCELL_82_808 ();
 FILLCELL_X32 FILLCELL_82_840 ();
 FILLCELL_X32 FILLCELL_82_872 ();
 FILLCELL_X32 FILLCELL_82_904 ();
 FILLCELL_X8 FILLCELL_82_936 ();
 FILLCELL_X32 FILLCELL_82_947 ();
 FILLCELL_X32 FILLCELL_82_979 ();
 FILLCELL_X32 FILLCELL_82_1011 ();
 FILLCELL_X32 FILLCELL_82_1043 ();
 FILLCELL_X32 FILLCELL_82_1075 ();
 FILLCELL_X32 FILLCELL_82_1107 ();
 FILLCELL_X32 FILLCELL_82_1139 ();
 FILLCELL_X32 FILLCELL_82_1171 ();
 FILLCELL_X32 FILLCELL_82_1203 ();
 FILLCELL_X32 FILLCELL_82_1235 ();
 FILLCELL_X32 FILLCELL_82_1267 ();
 FILLCELL_X32 FILLCELL_82_1299 ();
 FILLCELL_X32 FILLCELL_82_1331 ();
 FILLCELL_X32 FILLCELL_82_1363 ();
 FILLCELL_X32 FILLCELL_82_1395 ();
 FILLCELL_X32 FILLCELL_82_1427 ();
 FILLCELL_X32 FILLCELL_82_1459 ();
 FILLCELL_X32 FILLCELL_82_1491 ();
 FILLCELL_X32 FILLCELL_82_1523 ();
 FILLCELL_X32 FILLCELL_82_1555 ();
 FILLCELL_X32 FILLCELL_82_1587 ();
 FILLCELL_X32 FILLCELL_82_1619 ();
 FILLCELL_X32 FILLCELL_82_1651 ();
 FILLCELL_X32 FILLCELL_82_1683 ();
 FILLCELL_X32 FILLCELL_82_1715 ();
 FILLCELL_X32 FILLCELL_82_1747 ();
 FILLCELL_X32 FILLCELL_82_1779 ();
 FILLCELL_X32 FILLCELL_82_1811 ();
 FILLCELL_X32 FILLCELL_82_1843 ();
 FILLCELL_X16 FILLCELL_82_1875 ();
 FILLCELL_X4 FILLCELL_82_1891 ();
 FILLCELL_X2 FILLCELL_82_1895 ();
 FILLCELL_X32 FILLCELL_83_0 ();
 FILLCELL_X32 FILLCELL_83_32 ();
 FILLCELL_X32 FILLCELL_83_64 ();
 FILLCELL_X32 FILLCELL_83_96 ();
 FILLCELL_X32 FILLCELL_83_128 ();
 FILLCELL_X32 FILLCELL_83_160 ();
 FILLCELL_X32 FILLCELL_83_192 ();
 FILLCELL_X16 FILLCELL_83_224 ();
 FILLCELL_X4 FILLCELL_83_240 ();
 FILLCELL_X32 FILLCELL_83_247 ();
 FILLCELL_X32 FILLCELL_83_279 ();
 FILLCELL_X32 FILLCELL_83_311 ();
 FILLCELL_X32 FILLCELL_83_343 ();
 FILLCELL_X32 FILLCELL_83_375 ();
 FILLCELL_X32 FILLCELL_83_407 ();
 FILLCELL_X32 FILLCELL_83_439 ();
 FILLCELL_X32 FILLCELL_83_471 ();
 FILLCELL_X32 FILLCELL_83_503 ();
 FILLCELL_X32 FILLCELL_83_535 ();
 FILLCELL_X32 FILLCELL_83_567 ();
 FILLCELL_X32 FILLCELL_83_599 ();
 FILLCELL_X32 FILLCELL_83_631 ();
 FILLCELL_X32 FILLCELL_83_663 ();
 FILLCELL_X16 FILLCELL_83_695 ();
 FILLCELL_X8 FILLCELL_83_711 ();
 FILLCELL_X2 FILLCELL_83_719 ();
 FILLCELL_X32 FILLCELL_83_724 ();
 FILLCELL_X32 FILLCELL_83_756 ();
 FILLCELL_X32 FILLCELL_83_788 ();
 FILLCELL_X32 FILLCELL_83_820 ();
 FILLCELL_X32 FILLCELL_83_852 ();
 FILLCELL_X32 FILLCELL_83_884 ();
 FILLCELL_X32 FILLCELL_83_916 ();
 FILLCELL_X32 FILLCELL_83_948 ();
 FILLCELL_X32 FILLCELL_83_980 ();
 FILLCELL_X32 FILLCELL_83_1012 ();
 FILLCELL_X32 FILLCELL_83_1044 ();
 FILLCELL_X32 FILLCELL_83_1076 ();
 FILLCELL_X32 FILLCELL_83_1108 ();
 FILLCELL_X32 FILLCELL_83_1140 ();
 FILLCELL_X32 FILLCELL_83_1172 ();
 FILLCELL_X32 FILLCELL_83_1204 ();
 FILLCELL_X32 FILLCELL_83_1236 ();
 FILLCELL_X32 FILLCELL_83_1268 ();
 FILLCELL_X32 FILLCELL_83_1300 ();
 FILLCELL_X32 FILLCELL_83_1332 ();
 FILLCELL_X32 FILLCELL_83_1364 ();
 FILLCELL_X32 FILLCELL_83_1396 ();
 FILLCELL_X32 FILLCELL_83_1428 ();
 FILLCELL_X32 FILLCELL_83_1460 ();
 FILLCELL_X32 FILLCELL_83_1492 ();
 FILLCELL_X32 FILLCELL_83_1524 ();
 FILLCELL_X32 FILLCELL_83_1556 ();
 FILLCELL_X32 FILLCELL_83_1588 ();
 FILLCELL_X32 FILLCELL_83_1620 ();
 FILLCELL_X32 FILLCELL_83_1652 ();
 FILLCELL_X32 FILLCELL_83_1684 ();
 FILLCELL_X32 FILLCELL_83_1716 ();
 FILLCELL_X32 FILLCELL_83_1748 ();
 FILLCELL_X32 FILLCELL_83_1780 ();
 FILLCELL_X32 FILLCELL_83_1812 ();
 FILLCELL_X32 FILLCELL_83_1844 ();
 FILLCELL_X16 FILLCELL_83_1876 ();
 FILLCELL_X4 FILLCELL_83_1892 ();
 FILLCELL_X1 FILLCELL_83_1896 ();
 FILLCELL_X32 FILLCELL_84_0 ();
 FILLCELL_X32 FILLCELL_84_32 ();
 FILLCELL_X32 FILLCELL_84_64 ();
 FILLCELL_X32 FILLCELL_84_96 ();
 FILLCELL_X32 FILLCELL_84_128 ();
 FILLCELL_X32 FILLCELL_84_160 ();
 FILLCELL_X32 FILLCELL_84_192 ();
 FILLCELL_X32 FILLCELL_84_224 ();
 FILLCELL_X32 FILLCELL_84_256 ();
 FILLCELL_X32 FILLCELL_84_288 ();
 FILLCELL_X32 FILLCELL_84_320 ();
 FILLCELL_X32 FILLCELL_84_352 ();
 FILLCELL_X32 FILLCELL_84_384 ();
 FILLCELL_X32 FILLCELL_84_416 ();
 FILLCELL_X32 FILLCELL_84_448 ();
 FILLCELL_X32 FILLCELL_84_480 ();
 FILLCELL_X1 FILLCELL_84_512 ();
 FILLCELL_X32 FILLCELL_84_517 ();
 FILLCELL_X32 FILLCELL_84_549 ();
 FILLCELL_X32 FILLCELL_84_581 ();
 FILLCELL_X32 FILLCELL_84_613 ();
 FILLCELL_X32 FILLCELL_84_645 ();
 FILLCELL_X32 FILLCELL_84_677 ();
 FILLCELL_X32 FILLCELL_84_709 ();
 FILLCELL_X32 FILLCELL_84_741 ();
 FILLCELL_X32 FILLCELL_84_773 ();
 FILLCELL_X32 FILLCELL_84_805 ();
 FILLCELL_X32 FILLCELL_84_837 ();
 FILLCELL_X32 FILLCELL_84_869 ();
 FILLCELL_X32 FILLCELL_84_901 ();
 FILLCELL_X32 FILLCELL_84_933 ();
 FILLCELL_X32 FILLCELL_84_965 ();
 FILLCELL_X32 FILLCELL_84_997 ();
 FILLCELL_X32 FILLCELL_84_1029 ();
 FILLCELL_X32 FILLCELL_84_1061 ();
 FILLCELL_X32 FILLCELL_84_1093 ();
 FILLCELL_X32 FILLCELL_84_1125 ();
 FILLCELL_X32 FILLCELL_84_1157 ();
 FILLCELL_X32 FILLCELL_84_1189 ();
 FILLCELL_X32 FILLCELL_84_1221 ();
 FILLCELL_X32 FILLCELL_84_1253 ();
 FILLCELL_X32 FILLCELL_84_1285 ();
 FILLCELL_X32 FILLCELL_84_1317 ();
 FILLCELL_X32 FILLCELL_84_1349 ();
 FILLCELL_X32 FILLCELL_84_1381 ();
 FILLCELL_X32 FILLCELL_84_1413 ();
 FILLCELL_X32 FILLCELL_84_1445 ();
 FILLCELL_X32 FILLCELL_84_1477 ();
 FILLCELL_X32 FILLCELL_84_1509 ();
 FILLCELL_X32 FILLCELL_84_1541 ();
 FILLCELL_X32 FILLCELL_84_1573 ();
 FILLCELL_X32 FILLCELL_84_1605 ();
 FILLCELL_X32 FILLCELL_84_1637 ();
 FILLCELL_X32 FILLCELL_84_1669 ();
 FILLCELL_X32 FILLCELL_84_1701 ();
 FILLCELL_X32 FILLCELL_84_1733 ();
 FILLCELL_X32 FILLCELL_84_1765 ();
 FILLCELL_X32 FILLCELL_84_1797 ();
 FILLCELL_X32 FILLCELL_84_1829 ();
 FILLCELL_X32 FILLCELL_84_1861 ();
 FILLCELL_X4 FILLCELL_84_1893 ();
 FILLCELL_X32 FILLCELL_85_0 ();
 FILLCELL_X32 FILLCELL_85_32 ();
 FILLCELL_X32 FILLCELL_85_64 ();
 FILLCELL_X32 FILLCELL_85_96 ();
 FILLCELL_X32 FILLCELL_85_128 ();
 FILLCELL_X32 FILLCELL_85_160 ();
 FILLCELL_X32 FILLCELL_85_192 ();
 FILLCELL_X32 FILLCELL_85_224 ();
 FILLCELL_X32 FILLCELL_85_256 ();
 FILLCELL_X32 FILLCELL_85_288 ();
 FILLCELL_X32 FILLCELL_85_320 ();
 FILLCELL_X32 FILLCELL_85_352 ();
 FILLCELL_X32 FILLCELL_85_384 ();
 FILLCELL_X32 FILLCELL_85_416 ();
 FILLCELL_X32 FILLCELL_85_448 ();
 FILLCELL_X16 FILLCELL_85_480 ();
 FILLCELL_X4 FILLCELL_85_496 ();
 FILLCELL_X1 FILLCELL_85_500 ();
 FILLCELL_X32 FILLCELL_85_505 ();
 FILLCELL_X32 FILLCELL_85_537 ();
 FILLCELL_X32 FILLCELL_85_569 ();
 FILLCELL_X2 FILLCELL_85_601 ();
 FILLCELL_X1 FILLCELL_85_603 ();
 FILLCELL_X32 FILLCELL_85_607 ();
 FILLCELL_X32 FILLCELL_85_639 ();
 FILLCELL_X16 FILLCELL_85_671 ();
 FILLCELL_X32 FILLCELL_85_689 ();
 FILLCELL_X32 FILLCELL_85_721 ();
 FILLCELL_X32 FILLCELL_85_753 ();
 FILLCELL_X32 FILLCELL_85_785 ();
 FILLCELL_X16 FILLCELL_85_817 ();
 FILLCELL_X2 FILLCELL_85_833 ();
 FILLCELL_X1 FILLCELL_85_835 ();
 FILLCELL_X32 FILLCELL_85_853 ();
 FILLCELL_X32 FILLCELL_85_885 ();
 FILLCELL_X32 FILLCELL_85_917 ();
 FILLCELL_X32 FILLCELL_85_949 ();
 FILLCELL_X32 FILLCELL_85_981 ();
 FILLCELL_X32 FILLCELL_85_1013 ();
 FILLCELL_X32 FILLCELL_85_1045 ();
 FILLCELL_X32 FILLCELL_85_1077 ();
 FILLCELL_X32 FILLCELL_85_1109 ();
 FILLCELL_X32 FILLCELL_85_1141 ();
 FILLCELL_X32 FILLCELL_85_1173 ();
 FILLCELL_X32 FILLCELL_85_1205 ();
 FILLCELL_X32 FILLCELL_85_1237 ();
 FILLCELL_X32 FILLCELL_85_1269 ();
 FILLCELL_X32 FILLCELL_85_1301 ();
 FILLCELL_X32 FILLCELL_85_1333 ();
 FILLCELL_X32 FILLCELL_85_1365 ();
 FILLCELL_X32 FILLCELL_85_1397 ();
 FILLCELL_X32 FILLCELL_85_1429 ();
 FILLCELL_X32 FILLCELL_85_1461 ();
 FILLCELL_X32 FILLCELL_85_1493 ();
 FILLCELL_X32 FILLCELL_85_1525 ();
 FILLCELL_X32 FILLCELL_85_1557 ();
 FILLCELL_X32 FILLCELL_85_1589 ();
 FILLCELL_X32 FILLCELL_85_1621 ();
 FILLCELL_X32 FILLCELL_85_1653 ();
 FILLCELL_X32 FILLCELL_85_1685 ();
 FILLCELL_X32 FILLCELL_85_1717 ();
 FILLCELL_X32 FILLCELL_85_1749 ();
 FILLCELL_X32 FILLCELL_85_1781 ();
 FILLCELL_X32 FILLCELL_85_1813 ();
 FILLCELL_X32 FILLCELL_85_1845 ();
 FILLCELL_X16 FILLCELL_85_1877 ();
 FILLCELL_X4 FILLCELL_85_1893 ();
 FILLCELL_X32 FILLCELL_86_0 ();
 FILLCELL_X32 FILLCELL_86_32 ();
 FILLCELL_X32 FILLCELL_86_64 ();
 FILLCELL_X32 FILLCELL_86_96 ();
 FILLCELL_X32 FILLCELL_86_128 ();
 FILLCELL_X32 FILLCELL_86_160 ();
 FILLCELL_X32 FILLCELL_86_192 ();
 FILLCELL_X32 FILLCELL_86_224 ();
 FILLCELL_X32 FILLCELL_86_256 ();
 FILLCELL_X32 FILLCELL_86_288 ();
 FILLCELL_X32 FILLCELL_86_320 ();
 FILLCELL_X32 FILLCELL_86_352 ();
 FILLCELL_X32 FILLCELL_86_384 ();
 FILLCELL_X32 FILLCELL_86_416 ();
 FILLCELL_X32 FILLCELL_86_448 ();
 FILLCELL_X32 FILLCELL_86_480 ();
 FILLCELL_X32 FILLCELL_86_512 ();
 FILLCELL_X32 FILLCELL_86_544 ();
 FILLCELL_X32 FILLCELL_86_576 ();
 FILLCELL_X32 FILLCELL_86_608 ();
 FILLCELL_X32 FILLCELL_86_640 ();
 FILLCELL_X32 FILLCELL_86_672 ();
 FILLCELL_X32 FILLCELL_86_704 ();
 FILLCELL_X32 FILLCELL_86_736 ();
 FILLCELL_X32 FILLCELL_86_768 ();
 FILLCELL_X32 FILLCELL_86_800 ();
 FILLCELL_X32 FILLCELL_86_832 ();
 FILLCELL_X32 FILLCELL_86_864 ();
 FILLCELL_X32 FILLCELL_86_896 ();
 FILLCELL_X32 FILLCELL_86_928 ();
 FILLCELL_X32 FILLCELL_86_960 ();
 FILLCELL_X32 FILLCELL_86_992 ();
 FILLCELL_X32 FILLCELL_86_1024 ();
 FILLCELL_X32 FILLCELL_86_1056 ();
 FILLCELL_X32 FILLCELL_86_1088 ();
 FILLCELL_X32 FILLCELL_86_1120 ();
 FILLCELL_X32 FILLCELL_86_1152 ();
 FILLCELL_X32 FILLCELL_86_1184 ();
 FILLCELL_X32 FILLCELL_86_1216 ();
 FILLCELL_X32 FILLCELL_86_1248 ();
 FILLCELL_X32 FILLCELL_86_1280 ();
 FILLCELL_X32 FILLCELL_86_1312 ();
 FILLCELL_X32 FILLCELL_86_1344 ();
 FILLCELL_X32 FILLCELL_86_1376 ();
 FILLCELL_X32 FILLCELL_86_1408 ();
 FILLCELL_X32 FILLCELL_86_1440 ();
 FILLCELL_X32 FILLCELL_86_1472 ();
 FILLCELL_X32 FILLCELL_86_1504 ();
 FILLCELL_X32 FILLCELL_86_1536 ();
 FILLCELL_X32 FILLCELL_86_1568 ();
 FILLCELL_X32 FILLCELL_86_1600 ();
 FILLCELL_X32 FILLCELL_86_1632 ();
 FILLCELL_X32 FILLCELL_86_1664 ();
 FILLCELL_X32 FILLCELL_86_1696 ();
 FILLCELL_X32 FILLCELL_86_1728 ();
 FILLCELL_X32 FILLCELL_86_1760 ();
 FILLCELL_X32 FILLCELL_86_1792 ();
 FILLCELL_X32 FILLCELL_86_1824 ();
 FILLCELL_X32 FILLCELL_86_1856 ();
 FILLCELL_X8 FILLCELL_86_1888 ();
 FILLCELL_X1 FILLCELL_86_1896 ();
 FILLCELL_X32 FILLCELL_87_0 ();
 FILLCELL_X32 FILLCELL_87_32 ();
 FILLCELL_X32 FILLCELL_87_64 ();
 FILLCELL_X32 FILLCELL_87_96 ();
 FILLCELL_X32 FILLCELL_87_128 ();
 FILLCELL_X32 FILLCELL_87_160 ();
 FILLCELL_X32 FILLCELL_87_192 ();
 FILLCELL_X32 FILLCELL_87_224 ();
 FILLCELL_X32 FILLCELL_87_256 ();
 FILLCELL_X32 FILLCELL_87_288 ();
 FILLCELL_X32 FILLCELL_87_320 ();
 FILLCELL_X16 FILLCELL_87_352 ();
 FILLCELL_X8 FILLCELL_87_368 ();
 FILLCELL_X4 FILLCELL_87_376 ();
 FILLCELL_X2 FILLCELL_87_380 ();
 FILLCELL_X1 FILLCELL_87_382 ();
 FILLCELL_X32 FILLCELL_87_386 ();
 FILLCELL_X32 FILLCELL_87_418 ();
 FILLCELL_X32 FILLCELL_87_450 ();
 FILLCELL_X32 FILLCELL_87_482 ();
 FILLCELL_X32 FILLCELL_87_514 ();
 FILLCELL_X32 FILLCELL_87_546 ();
 FILLCELL_X32 FILLCELL_87_578 ();
 FILLCELL_X32 FILLCELL_87_610 ();
 FILLCELL_X32 FILLCELL_87_642 ();
 FILLCELL_X8 FILLCELL_87_674 ();
 FILLCELL_X4 FILLCELL_87_682 ();
 FILLCELL_X2 FILLCELL_87_686 ();
 FILLCELL_X32 FILLCELL_87_693 ();
 FILLCELL_X32 FILLCELL_87_725 ();
 FILLCELL_X32 FILLCELL_87_757 ();
 FILLCELL_X32 FILLCELL_87_789 ();
 FILLCELL_X32 FILLCELL_87_821 ();
 FILLCELL_X32 FILLCELL_87_853 ();
 FILLCELL_X32 FILLCELL_87_885 ();
 FILLCELL_X8 FILLCELL_87_917 ();
 FILLCELL_X2 FILLCELL_87_925 ();
 FILLCELL_X32 FILLCELL_87_930 ();
 FILLCELL_X32 FILLCELL_87_962 ();
 FILLCELL_X32 FILLCELL_87_994 ();
 FILLCELL_X32 FILLCELL_87_1026 ();
 FILLCELL_X32 FILLCELL_87_1058 ();
 FILLCELL_X32 FILLCELL_87_1090 ();
 FILLCELL_X32 FILLCELL_87_1122 ();
 FILLCELL_X32 FILLCELL_87_1154 ();
 FILLCELL_X32 FILLCELL_87_1186 ();
 FILLCELL_X32 FILLCELL_87_1218 ();
 FILLCELL_X32 FILLCELL_87_1250 ();
 FILLCELL_X32 FILLCELL_87_1282 ();
 FILLCELL_X32 FILLCELL_87_1314 ();
 FILLCELL_X32 FILLCELL_87_1346 ();
 FILLCELL_X32 FILLCELL_87_1378 ();
 FILLCELL_X32 FILLCELL_87_1410 ();
 FILLCELL_X32 FILLCELL_87_1442 ();
 FILLCELL_X32 FILLCELL_87_1474 ();
 FILLCELL_X32 FILLCELL_87_1506 ();
 FILLCELL_X32 FILLCELL_87_1538 ();
 FILLCELL_X32 FILLCELL_87_1570 ();
 FILLCELL_X32 FILLCELL_87_1602 ();
 FILLCELL_X32 FILLCELL_87_1634 ();
 FILLCELL_X32 FILLCELL_87_1666 ();
 FILLCELL_X32 FILLCELL_87_1698 ();
 FILLCELL_X32 FILLCELL_87_1730 ();
 FILLCELL_X32 FILLCELL_87_1762 ();
 FILLCELL_X32 FILLCELL_87_1794 ();
 FILLCELL_X32 FILLCELL_87_1826 ();
 FILLCELL_X32 FILLCELL_87_1858 ();
 FILLCELL_X4 FILLCELL_87_1890 ();
 FILLCELL_X2 FILLCELL_87_1894 ();
 FILLCELL_X1 FILLCELL_87_1896 ();
 FILLCELL_X32 FILLCELL_88_0 ();
 FILLCELL_X32 FILLCELL_88_32 ();
 FILLCELL_X32 FILLCELL_88_64 ();
 FILLCELL_X32 FILLCELL_88_96 ();
 FILLCELL_X32 FILLCELL_88_128 ();
 FILLCELL_X32 FILLCELL_88_160 ();
 FILLCELL_X32 FILLCELL_88_192 ();
 FILLCELL_X32 FILLCELL_88_224 ();
 FILLCELL_X32 FILLCELL_88_256 ();
 FILLCELL_X32 FILLCELL_88_288 ();
 FILLCELL_X32 FILLCELL_88_320 ();
 FILLCELL_X32 FILLCELL_88_352 ();
 FILLCELL_X32 FILLCELL_88_384 ();
 FILLCELL_X32 FILLCELL_88_416 ();
 FILLCELL_X32 FILLCELL_88_448 ();
 FILLCELL_X32 FILLCELL_88_480 ();
 FILLCELL_X8 FILLCELL_88_512 ();
 FILLCELL_X2 FILLCELL_88_520 ();
 FILLCELL_X32 FILLCELL_88_524 ();
 FILLCELL_X32 FILLCELL_88_556 ();
 FILLCELL_X32 FILLCELL_88_588 ();
 FILLCELL_X32 FILLCELL_88_620 ();
 FILLCELL_X32 FILLCELL_88_652 ();
 FILLCELL_X32 FILLCELL_88_684 ();
 FILLCELL_X32 FILLCELL_88_716 ();
 FILLCELL_X32 FILLCELL_88_748 ();
 FILLCELL_X32 FILLCELL_88_780 ();
 FILLCELL_X32 FILLCELL_88_812 ();
 FILLCELL_X32 FILLCELL_88_844 ();
 FILLCELL_X32 FILLCELL_88_876 ();
 FILLCELL_X32 FILLCELL_88_908 ();
 FILLCELL_X8 FILLCELL_88_940 ();
 FILLCELL_X4 FILLCELL_88_948 ();
 FILLCELL_X1 FILLCELL_88_952 ();
 FILLCELL_X32 FILLCELL_88_957 ();
 FILLCELL_X32 FILLCELL_88_989 ();
 FILLCELL_X32 FILLCELL_88_1021 ();
 FILLCELL_X32 FILLCELL_88_1053 ();
 FILLCELL_X32 FILLCELL_88_1085 ();
 FILLCELL_X32 FILLCELL_88_1117 ();
 FILLCELL_X32 FILLCELL_88_1149 ();
 FILLCELL_X32 FILLCELL_88_1181 ();
 FILLCELL_X32 FILLCELL_88_1213 ();
 FILLCELL_X32 FILLCELL_88_1245 ();
 FILLCELL_X32 FILLCELL_88_1277 ();
 FILLCELL_X32 FILLCELL_88_1309 ();
 FILLCELL_X32 FILLCELL_88_1341 ();
 FILLCELL_X32 FILLCELL_88_1373 ();
 FILLCELL_X32 FILLCELL_88_1405 ();
 FILLCELL_X32 FILLCELL_88_1437 ();
 FILLCELL_X32 FILLCELL_88_1469 ();
 FILLCELL_X32 FILLCELL_88_1501 ();
 FILLCELL_X32 FILLCELL_88_1533 ();
 FILLCELL_X32 FILLCELL_88_1565 ();
 FILLCELL_X32 FILLCELL_88_1597 ();
 FILLCELL_X32 FILLCELL_88_1629 ();
 FILLCELL_X32 FILLCELL_88_1661 ();
 FILLCELL_X32 FILLCELL_88_1693 ();
 FILLCELL_X32 FILLCELL_88_1725 ();
 FILLCELL_X32 FILLCELL_88_1757 ();
 FILLCELL_X32 FILLCELL_88_1789 ();
 FILLCELL_X32 FILLCELL_88_1821 ();
 FILLCELL_X32 FILLCELL_88_1853 ();
 FILLCELL_X8 FILLCELL_88_1885 ();
 FILLCELL_X4 FILLCELL_88_1893 ();
 FILLCELL_X32 FILLCELL_89_0 ();
 FILLCELL_X32 FILLCELL_89_32 ();
 FILLCELL_X32 FILLCELL_89_64 ();
 FILLCELL_X16 FILLCELL_89_96 ();
 FILLCELL_X8 FILLCELL_89_112 ();
 FILLCELL_X4 FILLCELL_89_120 ();
 FILLCELL_X2 FILLCELL_89_124 ();
 FILLCELL_X1 FILLCELL_89_126 ();
 FILLCELL_X32 FILLCELL_89_144 ();
 FILLCELL_X32 FILLCELL_89_176 ();
 FILLCELL_X32 FILLCELL_89_208 ();
 FILLCELL_X32 FILLCELL_89_240 ();
 FILLCELL_X32 FILLCELL_89_272 ();
 FILLCELL_X32 FILLCELL_89_304 ();
 FILLCELL_X32 FILLCELL_89_336 ();
 FILLCELL_X8 FILLCELL_89_368 ();
 FILLCELL_X4 FILLCELL_89_376 ();
 FILLCELL_X1 FILLCELL_89_380 ();
 FILLCELL_X32 FILLCELL_89_386 ();
 FILLCELL_X16 FILLCELL_89_418 ();
 FILLCELL_X2 FILLCELL_89_434 ();
 FILLCELL_X32 FILLCELL_89_438 ();
 FILLCELL_X32 FILLCELL_89_470 ();
 FILLCELL_X32 FILLCELL_89_502 ();
 FILLCELL_X32 FILLCELL_89_534 ();
 FILLCELL_X32 FILLCELL_89_566 ();
 FILLCELL_X32 FILLCELL_89_598 ();
 FILLCELL_X32 FILLCELL_89_630 ();
 FILLCELL_X4 FILLCELL_89_662 ();
 FILLCELL_X32 FILLCELL_89_670 ();
 FILLCELL_X32 FILLCELL_89_702 ();
 FILLCELL_X32 FILLCELL_89_734 ();
 FILLCELL_X32 FILLCELL_89_766 ();
 FILLCELL_X32 FILLCELL_89_798 ();
 FILLCELL_X2 FILLCELL_89_830 ();
 FILLCELL_X1 FILLCELL_89_832 ();
 FILLCELL_X32 FILLCELL_89_840 ();
 FILLCELL_X32 FILLCELL_89_872 ();
 FILLCELL_X32 FILLCELL_89_904 ();
 FILLCELL_X32 FILLCELL_89_936 ();
 FILLCELL_X32 FILLCELL_89_968 ();
 FILLCELL_X32 FILLCELL_89_1000 ();
 FILLCELL_X32 FILLCELL_89_1032 ();
 FILLCELL_X32 FILLCELL_89_1064 ();
 FILLCELL_X32 FILLCELL_89_1096 ();
 FILLCELL_X32 FILLCELL_89_1128 ();
 FILLCELL_X32 FILLCELL_89_1160 ();
 FILLCELL_X32 FILLCELL_89_1192 ();
 FILLCELL_X32 FILLCELL_89_1224 ();
 FILLCELL_X32 FILLCELL_89_1256 ();
 FILLCELL_X32 FILLCELL_89_1288 ();
 FILLCELL_X32 FILLCELL_89_1320 ();
 FILLCELL_X32 FILLCELL_89_1352 ();
 FILLCELL_X32 FILLCELL_89_1384 ();
 FILLCELL_X32 FILLCELL_89_1416 ();
 FILLCELL_X32 FILLCELL_89_1448 ();
 FILLCELL_X32 FILLCELL_89_1480 ();
 FILLCELL_X32 FILLCELL_89_1512 ();
 FILLCELL_X32 FILLCELL_89_1544 ();
 FILLCELL_X32 FILLCELL_89_1576 ();
 FILLCELL_X32 FILLCELL_89_1608 ();
 FILLCELL_X32 FILLCELL_89_1640 ();
 FILLCELL_X32 FILLCELL_89_1672 ();
 FILLCELL_X32 FILLCELL_89_1704 ();
 FILLCELL_X32 FILLCELL_89_1736 ();
 FILLCELL_X32 FILLCELL_89_1768 ();
 FILLCELL_X32 FILLCELL_89_1800 ();
 FILLCELL_X32 FILLCELL_89_1832 ();
 FILLCELL_X32 FILLCELL_89_1864 ();
 FILLCELL_X1 FILLCELL_89_1896 ();
 FILLCELL_X32 FILLCELL_90_0 ();
 FILLCELL_X32 FILLCELL_90_32 ();
 FILLCELL_X32 FILLCELL_90_64 ();
 FILLCELL_X32 FILLCELL_90_96 ();
 FILLCELL_X32 FILLCELL_90_128 ();
 FILLCELL_X16 FILLCELL_90_160 ();
 FILLCELL_X2 FILLCELL_90_176 ();
 FILLCELL_X4 FILLCELL_90_185 ();
 FILLCELL_X2 FILLCELL_90_189 ();
 FILLCELL_X1 FILLCELL_90_191 ();
 FILLCELL_X32 FILLCELL_90_194 ();
 FILLCELL_X32 FILLCELL_90_226 ();
 FILLCELL_X8 FILLCELL_90_258 ();
 FILLCELL_X2 FILLCELL_90_266 ();
 FILLCELL_X1 FILLCELL_90_268 ();
 FILLCELL_X8 FILLCELL_90_272 ();
 FILLCELL_X4 FILLCELL_90_280 ();
 FILLCELL_X2 FILLCELL_90_284 ();
 FILLCELL_X32 FILLCELL_90_289 ();
 FILLCELL_X8 FILLCELL_90_321 ();
 FILLCELL_X32 FILLCELL_90_333 ();
 FILLCELL_X16 FILLCELL_90_365 ();
 FILLCELL_X8 FILLCELL_90_381 ();
 FILLCELL_X4 FILLCELL_90_389 ();
 FILLCELL_X2 FILLCELL_90_393 ();
 FILLCELL_X32 FILLCELL_90_399 ();
 FILLCELL_X32 FILLCELL_90_431 ();
 FILLCELL_X32 FILLCELL_90_463 ();
 FILLCELL_X32 FILLCELL_90_495 ();
 FILLCELL_X32 FILLCELL_90_527 ();
 FILLCELL_X32 FILLCELL_90_559 ();
 FILLCELL_X32 FILLCELL_90_591 ();
 FILLCELL_X32 FILLCELL_90_623 ();
 FILLCELL_X32 FILLCELL_90_655 ();
 FILLCELL_X32 FILLCELL_90_687 ();
 FILLCELL_X16 FILLCELL_90_719 ();
 FILLCELL_X2 FILLCELL_90_735 ();
 FILLCELL_X32 FILLCELL_90_741 ();
 FILLCELL_X32 FILLCELL_90_773 ();
 FILLCELL_X32 FILLCELL_90_805 ();
 FILLCELL_X32 FILLCELL_90_837 ();
 FILLCELL_X32 FILLCELL_90_869 ();
 FILLCELL_X32 FILLCELL_90_901 ();
 FILLCELL_X16 FILLCELL_90_933 ();
 FILLCELL_X8 FILLCELL_90_949 ();
 FILLCELL_X4 FILLCELL_90_957 ();
 FILLCELL_X2 FILLCELL_90_961 ();
 FILLCELL_X32 FILLCELL_90_968 ();
 FILLCELL_X32 FILLCELL_90_1000 ();
 FILLCELL_X32 FILLCELL_90_1032 ();
 FILLCELL_X32 FILLCELL_90_1064 ();
 FILLCELL_X32 FILLCELL_90_1096 ();
 FILLCELL_X32 FILLCELL_90_1128 ();
 FILLCELL_X32 FILLCELL_90_1160 ();
 FILLCELL_X32 FILLCELL_90_1192 ();
 FILLCELL_X32 FILLCELL_90_1224 ();
 FILLCELL_X32 FILLCELL_90_1256 ();
 FILLCELL_X32 FILLCELL_90_1288 ();
 FILLCELL_X32 FILLCELL_90_1320 ();
 FILLCELL_X32 FILLCELL_90_1352 ();
 FILLCELL_X32 FILLCELL_90_1384 ();
 FILLCELL_X32 FILLCELL_90_1416 ();
 FILLCELL_X32 FILLCELL_90_1448 ();
 FILLCELL_X32 FILLCELL_90_1480 ();
 FILLCELL_X32 FILLCELL_90_1512 ();
 FILLCELL_X32 FILLCELL_90_1544 ();
 FILLCELL_X32 FILLCELL_90_1576 ();
 FILLCELL_X32 FILLCELL_90_1608 ();
 FILLCELL_X32 FILLCELL_90_1640 ();
 FILLCELL_X32 FILLCELL_90_1672 ();
 FILLCELL_X32 FILLCELL_90_1704 ();
 FILLCELL_X32 FILLCELL_90_1736 ();
 FILLCELL_X32 FILLCELL_90_1768 ();
 FILLCELL_X32 FILLCELL_90_1800 ();
 FILLCELL_X32 FILLCELL_90_1832 ();
 FILLCELL_X32 FILLCELL_90_1864 ();
 FILLCELL_X1 FILLCELL_90_1896 ();
 FILLCELL_X32 FILLCELL_91_0 ();
 FILLCELL_X32 FILLCELL_91_32 ();
 FILLCELL_X32 FILLCELL_91_64 ();
 FILLCELL_X32 FILLCELL_91_96 ();
 FILLCELL_X32 FILLCELL_91_128 ();
 FILLCELL_X32 FILLCELL_91_160 ();
 FILLCELL_X32 FILLCELL_91_192 ();
 FILLCELL_X32 FILLCELL_91_224 ();
 FILLCELL_X32 FILLCELL_91_256 ();
 FILLCELL_X32 FILLCELL_91_288 ();
 FILLCELL_X16 FILLCELL_91_320 ();
 FILLCELL_X8 FILLCELL_91_336 ();
 FILLCELL_X4 FILLCELL_91_344 ();
 FILLCELL_X1 FILLCELL_91_348 ();
 FILLCELL_X32 FILLCELL_91_351 ();
 FILLCELL_X32 FILLCELL_91_383 ();
 FILLCELL_X32 FILLCELL_91_415 ();
 FILLCELL_X32 FILLCELL_91_447 ();
 FILLCELL_X16 FILLCELL_91_479 ();
 FILLCELL_X8 FILLCELL_91_495 ();
 FILLCELL_X4 FILLCELL_91_503 ();
 FILLCELL_X2 FILLCELL_91_507 ();
 FILLCELL_X32 FILLCELL_91_513 ();
 FILLCELL_X32 FILLCELL_91_545 ();
 FILLCELL_X32 FILLCELL_91_577 ();
 FILLCELL_X32 FILLCELL_91_609 ();
 FILLCELL_X32 FILLCELL_91_641 ();
 FILLCELL_X32 FILLCELL_91_673 ();
 FILLCELL_X32 FILLCELL_91_705 ();
 FILLCELL_X32 FILLCELL_91_737 ();
 FILLCELL_X32 FILLCELL_91_769 ();
 FILLCELL_X32 FILLCELL_91_801 ();
 FILLCELL_X32 FILLCELL_91_833 ();
 FILLCELL_X32 FILLCELL_91_865 ();
 FILLCELL_X32 FILLCELL_91_897 ();
 FILLCELL_X16 FILLCELL_91_929 ();
 FILLCELL_X4 FILLCELL_91_945 ();
 FILLCELL_X2 FILLCELL_91_949 ();
 FILLCELL_X32 FILLCELL_91_953 ();
 FILLCELL_X32 FILLCELL_91_985 ();
 FILLCELL_X32 FILLCELL_91_1017 ();
 FILLCELL_X32 FILLCELL_91_1049 ();
 FILLCELL_X32 FILLCELL_91_1081 ();
 FILLCELL_X32 FILLCELL_91_1113 ();
 FILLCELL_X32 FILLCELL_91_1145 ();
 FILLCELL_X32 FILLCELL_91_1177 ();
 FILLCELL_X32 FILLCELL_91_1209 ();
 FILLCELL_X32 FILLCELL_91_1241 ();
 FILLCELL_X32 FILLCELL_91_1273 ();
 FILLCELL_X32 FILLCELL_91_1305 ();
 FILLCELL_X32 FILLCELL_91_1337 ();
 FILLCELL_X32 FILLCELL_91_1369 ();
 FILLCELL_X32 FILLCELL_91_1401 ();
 FILLCELL_X32 FILLCELL_91_1433 ();
 FILLCELL_X32 FILLCELL_91_1465 ();
 FILLCELL_X32 FILLCELL_91_1497 ();
 FILLCELL_X32 FILLCELL_91_1529 ();
 FILLCELL_X32 FILLCELL_91_1561 ();
 FILLCELL_X32 FILLCELL_91_1593 ();
 FILLCELL_X32 FILLCELL_91_1625 ();
 FILLCELL_X32 FILLCELL_91_1657 ();
 FILLCELL_X32 FILLCELL_91_1689 ();
 FILLCELL_X32 FILLCELL_91_1721 ();
 FILLCELL_X32 FILLCELL_91_1753 ();
 FILLCELL_X32 FILLCELL_91_1785 ();
 FILLCELL_X32 FILLCELL_91_1817 ();
 FILLCELL_X32 FILLCELL_91_1849 ();
 FILLCELL_X16 FILLCELL_91_1881 ();
 FILLCELL_X32 FILLCELL_92_0 ();
 FILLCELL_X32 FILLCELL_92_32 ();
 FILLCELL_X32 FILLCELL_92_64 ();
 FILLCELL_X32 FILLCELL_92_96 ();
 FILLCELL_X32 FILLCELL_92_128 ();
 FILLCELL_X32 FILLCELL_92_160 ();
 FILLCELL_X32 FILLCELL_92_192 ();
 FILLCELL_X32 FILLCELL_92_224 ();
 FILLCELL_X32 FILLCELL_92_256 ();
 FILLCELL_X32 FILLCELL_92_288 ();
 FILLCELL_X32 FILLCELL_92_320 ();
 FILLCELL_X32 FILLCELL_92_352 ();
 FILLCELL_X32 FILLCELL_92_384 ();
 FILLCELL_X32 FILLCELL_92_416 ();
 FILLCELL_X32 FILLCELL_92_448 ();
 FILLCELL_X32 FILLCELL_92_480 ();
 FILLCELL_X32 FILLCELL_92_512 ();
 FILLCELL_X32 FILLCELL_92_544 ();
 FILLCELL_X32 FILLCELL_92_576 ();
 FILLCELL_X32 FILLCELL_92_608 ();
 FILLCELL_X32 FILLCELL_92_640 ();
 FILLCELL_X32 FILLCELL_92_672 ();
 FILLCELL_X32 FILLCELL_92_704 ();
 FILLCELL_X32 FILLCELL_92_741 ();
 FILLCELL_X32 FILLCELL_92_773 ();
 FILLCELL_X16 FILLCELL_92_805 ();
 FILLCELL_X4 FILLCELL_92_821 ();
 FILLCELL_X16 FILLCELL_92_830 ();
 FILLCELL_X4 FILLCELL_92_846 ();
 FILLCELL_X2 FILLCELL_92_850 ();
 FILLCELL_X32 FILLCELL_92_855 ();
 FILLCELL_X32 FILLCELL_92_887 ();
 FILLCELL_X32 FILLCELL_92_919 ();
 FILLCELL_X32 FILLCELL_92_951 ();
 FILLCELL_X32 FILLCELL_92_983 ();
 FILLCELL_X32 FILLCELL_92_1015 ();
 FILLCELL_X32 FILLCELL_92_1047 ();
 FILLCELL_X32 FILLCELL_92_1079 ();
 FILLCELL_X32 FILLCELL_92_1111 ();
 FILLCELL_X32 FILLCELL_92_1143 ();
 FILLCELL_X32 FILLCELL_92_1175 ();
 FILLCELL_X32 FILLCELL_92_1207 ();
 FILLCELL_X32 FILLCELL_92_1239 ();
 FILLCELL_X32 FILLCELL_92_1271 ();
 FILLCELL_X32 FILLCELL_92_1303 ();
 FILLCELL_X32 FILLCELL_92_1335 ();
 FILLCELL_X32 FILLCELL_92_1367 ();
 FILLCELL_X32 FILLCELL_92_1399 ();
 FILLCELL_X32 FILLCELL_92_1431 ();
 FILLCELL_X32 FILLCELL_92_1463 ();
 FILLCELL_X32 FILLCELL_92_1495 ();
 FILLCELL_X32 FILLCELL_92_1527 ();
 FILLCELL_X32 FILLCELL_92_1559 ();
 FILLCELL_X32 FILLCELL_92_1591 ();
 FILLCELL_X32 FILLCELL_92_1623 ();
 FILLCELL_X32 FILLCELL_92_1655 ();
 FILLCELL_X32 FILLCELL_92_1687 ();
 FILLCELL_X32 FILLCELL_92_1719 ();
 FILLCELL_X32 FILLCELL_92_1751 ();
 FILLCELL_X32 FILLCELL_92_1783 ();
 FILLCELL_X32 FILLCELL_92_1815 ();
 FILLCELL_X32 FILLCELL_92_1847 ();
 FILLCELL_X16 FILLCELL_92_1879 ();
 FILLCELL_X2 FILLCELL_92_1895 ();
 FILLCELL_X32 FILLCELL_93_0 ();
 FILLCELL_X32 FILLCELL_93_32 ();
 FILLCELL_X32 FILLCELL_93_64 ();
 FILLCELL_X32 FILLCELL_93_96 ();
 FILLCELL_X32 FILLCELL_93_128 ();
 FILLCELL_X32 FILLCELL_93_160 ();
 FILLCELL_X32 FILLCELL_93_192 ();
 FILLCELL_X16 FILLCELL_93_224 ();
 FILLCELL_X2 FILLCELL_93_240 ();
 FILLCELL_X1 FILLCELL_93_242 ();
 FILLCELL_X4 FILLCELL_93_247 ();
 FILLCELL_X32 FILLCELL_93_257 ();
 FILLCELL_X32 FILLCELL_93_289 ();
 FILLCELL_X32 FILLCELL_93_321 ();
 FILLCELL_X32 FILLCELL_93_353 ();
 FILLCELL_X8 FILLCELL_93_385 ();
 FILLCELL_X2 FILLCELL_93_393 ();
 FILLCELL_X32 FILLCELL_93_398 ();
 FILLCELL_X32 FILLCELL_93_430 ();
 FILLCELL_X32 FILLCELL_93_462 ();
 FILLCELL_X32 FILLCELL_93_494 ();
 FILLCELL_X32 FILLCELL_93_526 ();
 FILLCELL_X32 FILLCELL_93_558 ();
 FILLCELL_X32 FILLCELL_93_590 ();
 FILLCELL_X16 FILLCELL_93_622 ();
 FILLCELL_X8 FILLCELL_93_638 ();
 FILLCELL_X32 FILLCELL_93_649 ();
 FILLCELL_X32 FILLCELL_93_681 ();
 FILLCELL_X32 FILLCELL_93_713 ();
 FILLCELL_X32 FILLCELL_93_745 ();
 FILLCELL_X32 FILLCELL_93_777 ();
 FILLCELL_X32 FILLCELL_93_809 ();
 FILLCELL_X2 FILLCELL_93_841 ();
 FILLCELL_X32 FILLCELL_93_849 ();
 FILLCELL_X32 FILLCELL_93_881 ();
 FILLCELL_X32 FILLCELL_93_913 ();
 FILLCELL_X32 FILLCELL_93_945 ();
 FILLCELL_X32 FILLCELL_93_977 ();
 FILLCELL_X32 FILLCELL_93_1009 ();
 FILLCELL_X32 FILLCELL_93_1041 ();
 FILLCELL_X32 FILLCELL_93_1073 ();
 FILLCELL_X32 FILLCELL_93_1105 ();
 FILLCELL_X32 FILLCELL_93_1137 ();
 FILLCELL_X32 FILLCELL_93_1169 ();
 FILLCELL_X32 FILLCELL_93_1201 ();
 FILLCELL_X32 FILLCELL_93_1233 ();
 FILLCELL_X32 FILLCELL_93_1265 ();
 FILLCELL_X32 FILLCELL_93_1297 ();
 FILLCELL_X32 FILLCELL_93_1329 ();
 FILLCELL_X32 FILLCELL_93_1361 ();
 FILLCELL_X32 FILLCELL_93_1393 ();
 FILLCELL_X32 FILLCELL_93_1425 ();
 FILLCELL_X32 FILLCELL_93_1457 ();
 FILLCELL_X32 FILLCELL_93_1489 ();
 FILLCELL_X32 FILLCELL_93_1521 ();
 FILLCELL_X32 FILLCELL_93_1553 ();
 FILLCELL_X32 FILLCELL_93_1585 ();
 FILLCELL_X32 FILLCELL_93_1617 ();
 FILLCELL_X32 FILLCELL_93_1649 ();
 FILLCELL_X32 FILLCELL_93_1681 ();
 FILLCELL_X32 FILLCELL_93_1713 ();
 FILLCELL_X32 FILLCELL_93_1745 ();
 FILLCELL_X32 FILLCELL_93_1777 ();
 FILLCELL_X32 FILLCELL_93_1809 ();
 FILLCELL_X32 FILLCELL_93_1841 ();
 FILLCELL_X16 FILLCELL_93_1873 ();
 FILLCELL_X8 FILLCELL_93_1889 ();
 FILLCELL_X32 FILLCELL_94_0 ();
 FILLCELL_X32 FILLCELL_94_32 ();
 FILLCELL_X32 FILLCELL_94_64 ();
 FILLCELL_X32 FILLCELL_94_96 ();
 FILLCELL_X32 FILLCELL_94_128 ();
 FILLCELL_X32 FILLCELL_94_160 ();
 FILLCELL_X32 FILLCELL_94_192 ();
 FILLCELL_X16 FILLCELL_94_224 ();
 FILLCELL_X32 FILLCELL_94_243 ();
 FILLCELL_X32 FILLCELL_94_275 ();
 FILLCELL_X32 FILLCELL_94_307 ();
 FILLCELL_X32 FILLCELL_94_339 ();
 FILLCELL_X32 FILLCELL_94_371 ();
 FILLCELL_X32 FILLCELL_94_403 ();
 FILLCELL_X32 FILLCELL_94_435 ();
 FILLCELL_X32 FILLCELL_94_467 ();
 FILLCELL_X16 FILLCELL_94_499 ();
 FILLCELL_X1 FILLCELL_94_515 ();
 FILLCELL_X32 FILLCELL_94_519 ();
 FILLCELL_X32 FILLCELL_94_551 ();
 FILLCELL_X32 FILLCELL_94_583 ();
 FILLCELL_X16 FILLCELL_94_615 ();
 FILLCELL_X4 FILLCELL_94_631 ();
 FILLCELL_X32 FILLCELL_94_637 ();
 FILLCELL_X32 FILLCELL_94_669 ();
 FILLCELL_X32 FILLCELL_94_701 ();
 FILLCELL_X32 FILLCELL_94_733 ();
 FILLCELL_X32 FILLCELL_94_765 ();
 FILLCELL_X32 FILLCELL_94_797 ();
 FILLCELL_X32 FILLCELL_94_829 ();
 FILLCELL_X32 FILLCELL_94_861 ();
 FILLCELL_X32 FILLCELL_94_893 ();
 FILLCELL_X32 FILLCELL_94_925 ();
 FILLCELL_X32 FILLCELL_94_957 ();
 FILLCELL_X32 FILLCELL_94_989 ();
 FILLCELL_X32 FILLCELL_94_1021 ();
 FILLCELL_X32 FILLCELL_94_1053 ();
 FILLCELL_X32 FILLCELL_94_1085 ();
 FILLCELL_X32 FILLCELL_94_1117 ();
 FILLCELL_X32 FILLCELL_94_1149 ();
 FILLCELL_X32 FILLCELL_94_1181 ();
 FILLCELL_X32 FILLCELL_94_1213 ();
 FILLCELL_X32 FILLCELL_94_1245 ();
 FILLCELL_X32 FILLCELL_94_1277 ();
 FILLCELL_X32 FILLCELL_94_1309 ();
 FILLCELL_X32 FILLCELL_94_1341 ();
 FILLCELL_X32 FILLCELL_94_1373 ();
 FILLCELL_X32 FILLCELL_94_1405 ();
 FILLCELL_X32 FILLCELL_94_1437 ();
 FILLCELL_X32 FILLCELL_94_1469 ();
 FILLCELL_X32 FILLCELL_94_1501 ();
 FILLCELL_X32 FILLCELL_94_1533 ();
 FILLCELL_X32 FILLCELL_94_1565 ();
 FILLCELL_X32 FILLCELL_94_1597 ();
 FILLCELL_X32 FILLCELL_94_1629 ();
 FILLCELL_X32 FILLCELL_94_1661 ();
 FILLCELL_X32 FILLCELL_94_1693 ();
 FILLCELL_X32 FILLCELL_94_1725 ();
 FILLCELL_X32 FILLCELL_94_1757 ();
 FILLCELL_X32 FILLCELL_94_1789 ();
 FILLCELL_X32 FILLCELL_94_1821 ();
 FILLCELL_X32 FILLCELL_94_1853 ();
 FILLCELL_X8 FILLCELL_94_1885 ();
 FILLCELL_X4 FILLCELL_94_1893 ();
 FILLCELL_X32 FILLCELL_95_0 ();
 FILLCELL_X32 FILLCELL_95_32 ();
 FILLCELL_X32 FILLCELL_95_64 ();
 FILLCELL_X32 FILLCELL_95_96 ();
 FILLCELL_X32 FILLCELL_95_128 ();
 FILLCELL_X32 FILLCELL_95_160 ();
 FILLCELL_X32 FILLCELL_95_192 ();
 FILLCELL_X32 FILLCELL_95_224 ();
 FILLCELL_X32 FILLCELL_95_256 ();
 FILLCELL_X32 FILLCELL_95_288 ();
 FILLCELL_X4 FILLCELL_95_320 ();
 FILLCELL_X2 FILLCELL_95_324 ();
 FILLCELL_X1 FILLCELL_95_326 ();
 FILLCELL_X32 FILLCELL_95_330 ();
 FILLCELL_X32 FILLCELL_95_362 ();
 FILLCELL_X32 FILLCELL_95_394 ();
 FILLCELL_X32 FILLCELL_95_426 ();
 FILLCELL_X32 FILLCELL_95_458 ();
 FILLCELL_X8 FILLCELL_95_490 ();
 FILLCELL_X2 FILLCELL_95_498 ();
 FILLCELL_X1 FILLCELL_95_500 ();
 FILLCELL_X32 FILLCELL_95_504 ();
 FILLCELL_X32 FILLCELL_95_536 ();
 FILLCELL_X32 FILLCELL_95_568 ();
 FILLCELL_X16 FILLCELL_95_600 ();
 FILLCELL_X4 FILLCELL_95_616 ();
 FILLCELL_X2 FILLCELL_95_620 ();
 FILLCELL_X16 FILLCELL_95_625 ();
 FILLCELL_X8 FILLCELL_95_641 ();
 FILLCELL_X4 FILLCELL_95_649 ();
 FILLCELL_X2 FILLCELL_95_653 ();
 FILLCELL_X1 FILLCELL_95_655 ();
 FILLCELL_X32 FILLCELL_95_659 ();
 FILLCELL_X32 FILLCELL_95_691 ();
 FILLCELL_X32 FILLCELL_95_723 ();
 FILLCELL_X32 FILLCELL_95_755 ();
 FILLCELL_X32 FILLCELL_95_787 ();
 FILLCELL_X32 FILLCELL_95_819 ();
 FILLCELL_X32 FILLCELL_95_851 ();
 FILLCELL_X32 FILLCELL_95_883 ();
 FILLCELL_X32 FILLCELL_95_915 ();
 FILLCELL_X32 FILLCELL_95_947 ();
 FILLCELL_X1 FILLCELL_95_979 ();
 FILLCELL_X32 FILLCELL_95_987 ();
 FILLCELL_X32 FILLCELL_95_1019 ();
 FILLCELL_X32 FILLCELL_95_1051 ();
 FILLCELL_X32 FILLCELL_95_1083 ();
 FILLCELL_X32 FILLCELL_95_1115 ();
 FILLCELL_X32 FILLCELL_95_1147 ();
 FILLCELL_X32 FILLCELL_95_1179 ();
 FILLCELL_X32 FILLCELL_95_1211 ();
 FILLCELL_X32 FILLCELL_95_1243 ();
 FILLCELL_X32 FILLCELL_95_1275 ();
 FILLCELL_X32 FILLCELL_95_1307 ();
 FILLCELL_X32 FILLCELL_95_1339 ();
 FILLCELL_X32 FILLCELL_95_1371 ();
 FILLCELL_X32 FILLCELL_95_1403 ();
 FILLCELL_X32 FILLCELL_95_1435 ();
 FILLCELL_X32 FILLCELL_95_1467 ();
 FILLCELL_X32 FILLCELL_95_1499 ();
 FILLCELL_X32 FILLCELL_95_1531 ();
 FILLCELL_X32 FILLCELL_95_1563 ();
 FILLCELL_X32 FILLCELL_95_1595 ();
 FILLCELL_X32 FILLCELL_95_1627 ();
 FILLCELL_X32 FILLCELL_95_1659 ();
 FILLCELL_X32 FILLCELL_95_1691 ();
 FILLCELL_X32 FILLCELL_95_1723 ();
 FILLCELL_X32 FILLCELL_95_1755 ();
 FILLCELL_X32 FILLCELL_95_1787 ();
 FILLCELL_X32 FILLCELL_95_1819 ();
 FILLCELL_X32 FILLCELL_95_1851 ();
 FILLCELL_X8 FILLCELL_95_1883 ();
 FILLCELL_X4 FILLCELL_95_1891 ();
 FILLCELL_X2 FILLCELL_95_1895 ();
 FILLCELL_X32 FILLCELL_96_0 ();
 FILLCELL_X32 FILLCELL_96_32 ();
 FILLCELL_X32 FILLCELL_96_64 ();
 FILLCELL_X32 FILLCELL_96_96 ();
 FILLCELL_X32 FILLCELL_96_128 ();
 FILLCELL_X32 FILLCELL_96_160 ();
 FILLCELL_X32 FILLCELL_96_192 ();
 FILLCELL_X32 FILLCELL_96_224 ();
 FILLCELL_X32 FILLCELL_96_256 ();
 FILLCELL_X32 FILLCELL_96_288 ();
 FILLCELL_X32 FILLCELL_96_320 ();
 FILLCELL_X2 FILLCELL_96_352 ();
 FILLCELL_X1 FILLCELL_96_354 ();
 FILLCELL_X32 FILLCELL_96_358 ();
 FILLCELL_X32 FILLCELL_96_390 ();
 FILLCELL_X32 FILLCELL_96_422 ();
 FILLCELL_X32 FILLCELL_96_454 ();
 FILLCELL_X32 FILLCELL_96_486 ();
 FILLCELL_X32 FILLCELL_96_518 ();
 FILLCELL_X32 FILLCELL_96_550 ();
 FILLCELL_X32 FILLCELL_96_582 ();
 FILLCELL_X32 FILLCELL_96_614 ();
 FILLCELL_X32 FILLCELL_96_646 ();
 FILLCELL_X32 FILLCELL_96_678 ();
 FILLCELL_X32 FILLCELL_96_710 ();
 FILLCELL_X32 FILLCELL_96_742 ();
 FILLCELL_X32 FILLCELL_96_774 ();
 FILLCELL_X32 FILLCELL_96_806 ();
 FILLCELL_X32 FILLCELL_96_838 ();
 FILLCELL_X32 FILLCELL_96_870 ();
 FILLCELL_X32 FILLCELL_96_902 ();
 FILLCELL_X32 FILLCELL_96_934 ();
 FILLCELL_X32 FILLCELL_96_966 ();
 FILLCELL_X32 FILLCELL_96_998 ();
 FILLCELL_X8 FILLCELL_96_1030 ();
 FILLCELL_X4 FILLCELL_96_1038 ();
 FILLCELL_X2 FILLCELL_96_1042 ();
 FILLCELL_X32 FILLCELL_96_1061 ();
 FILLCELL_X32 FILLCELL_96_1093 ();
 FILLCELL_X32 FILLCELL_96_1125 ();
 FILLCELL_X32 FILLCELL_96_1157 ();
 FILLCELL_X32 FILLCELL_96_1189 ();
 FILLCELL_X32 FILLCELL_96_1221 ();
 FILLCELL_X32 FILLCELL_96_1253 ();
 FILLCELL_X32 FILLCELL_96_1285 ();
 FILLCELL_X32 FILLCELL_96_1317 ();
 FILLCELL_X32 FILLCELL_96_1349 ();
 FILLCELL_X32 FILLCELL_96_1381 ();
 FILLCELL_X32 FILLCELL_96_1413 ();
 FILLCELL_X32 FILLCELL_96_1445 ();
 FILLCELL_X32 FILLCELL_96_1477 ();
 FILLCELL_X32 FILLCELL_96_1509 ();
 FILLCELL_X32 FILLCELL_96_1541 ();
 FILLCELL_X32 FILLCELL_96_1573 ();
 FILLCELL_X32 FILLCELL_96_1605 ();
 FILLCELL_X32 FILLCELL_96_1637 ();
 FILLCELL_X32 FILLCELL_96_1669 ();
 FILLCELL_X32 FILLCELL_96_1701 ();
 FILLCELL_X32 FILLCELL_96_1733 ();
 FILLCELL_X32 FILLCELL_96_1765 ();
 FILLCELL_X32 FILLCELL_96_1797 ();
 FILLCELL_X32 FILLCELL_96_1829 ();
 FILLCELL_X32 FILLCELL_96_1861 ();
 FILLCELL_X4 FILLCELL_96_1893 ();
 FILLCELL_X32 FILLCELL_97_0 ();
 FILLCELL_X32 FILLCELL_97_32 ();
 FILLCELL_X32 FILLCELL_97_64 ();
 FILLCELL_X32 FILLCELL_97_96 ();
 FILLCELL_X32 FILLCELL_97_128 ();
 FILLCELL_X32 FILLCELL_97_160 ();
 FILLCELL_X32 FILLCELL_97_192 ();
 FILLCELL_X32 FILLCELL_97_224 ();
 FILLCELL_X32 FILLCELL_97_256 ();
 FILLCELL_X32 FILLCELL_97_288 ();
 FILLCELL_X32 FILLCELL_97_320 ();
 FILLCELL_X32 FILLCELL_97_352 ();
 FILLCELL_X32 FILLCELL_97_384 ();
 FILLCELL_X32 FILLCELL_97_416 ();
 FILLCELL_X32 FILLCELL_97_448 ();
 FILLCELL_X32 FILLCELL_97_480 ();
 FILLCELL_X16 FILLCELL_97_512 ();
 FILLCELL_X8 FILLCELL_97_528 ();
 FILLCELL_X4 FILLCELL_97_536 ();
 FILLCELL_X2 FILLCELL_97_540 ();
 FILLCELL_X1 FILLCELL_97_542 ();
 FILLCELL_X8 FILLCELL_97_546 ();
 FILLCELL_X4 FILLCELL_97_554 ();
 FILLCELL_X2 FILLCELL_97_558 ();
 FILLCELL_X32 FILLCELL_97_563 ();
 FILLCELL_X32 FILLCELL_97_595 ();
 FILLCELL_X16 FILLCELL_97_627 ();
 FILLCELL_X2 FILLCELL_97_643 ();
 FILLCELL_X32 FILLCELL_97_649 ();
 FILLCELL_X32 FILLCELL_97_681 ();
 FILLCELL_X32 FILLCELL_97_713 ();
 FILLCELL_X32 FILLCELL_97_745 ();
 FILLCELL_X32 FILLCELL_97_777 ();
 FILLCELL_X8 FILLCELL_97_809 ();
 FILLCELL_X4 FILLCELL_97_817 ();
 FILLCELL_X1 FILLCELL_97_821 ();
 FILLCELL_X32 FILLCELL_97_826 ();
 FILLCELL_X32 FILLCELL_97_858 ();
 FILLCELL_X32 FILLCELL_97_890 ();
 FILLCELL_X32 FILLCELL_97_922 ();
 FILLCELL_X4 FILLCELL_97_954 ();
 FILLCELL_X2 FILLCELL_97_958 ();
 FILLCELL_X32 FILLCELL_97_963 ();
 FILLCELL_X32 FILLCELL_97_995 ();
 FILLCELL_X32 FILLCELL_97_1027 ();
 FILLCELL_X32 FILLCELL_97_1059 ();
 FILLCELL_X32 FILLCELL_97_1091 ();
 FILLCELL_X32 FILLCELL_97_1123 ();
 FILLCELL_X32 FILLCELL_97_1155 ();
 FILLCELL_X32 FILLCELL_97_1187 ();
 FILLCELL_X32 FILLCELL_97_1219 ();
 FILLCELL_X32 FILLCELL_97_1251 ();
 FILLCELL_X32 FILLCELL_97_1283 ();
 FILLCELL_X32 FILLCELL_97_1315 ();
 FILLCELL_X32 FILLCELL_97_1347 ();
 FILLCELL_X32 FILLCELL_97_1379 ();
 FILLCELL_X32 FILLCELL_97_1411 ();
 FILLCELL_X32 FILLCELL_97_1443 ();
 FILLCELL_X32 FILLCELL_97_1475 ();
 FILLCELL_X32 FILLCELL_97_1507 ();
 FILLCELL_X32 FILLCELL_97_1539 ();
 FILLCELL_X32 FILLCELL_97_1571 ();
 FILLCELL_X32 FILLCELL_97_1603 ();
 FILLCELL_X32 FILLCELL_97_1635 ();
 FILLCELL_X32 FILLCELL_97_1667 ();
 FILLCELL_X32 FILLCELL_97_1699 ();
 FILLCELL_X32 FILLCELL_97_1731 ();
 FILLCELL_X32 FILLCELL_97_1763 ();
 FILLCELL_X32 FILLCELL_97_1795 ();
 FILLCELL_X32 FILLCELL_97_1827 ();
 FILLCELL_X32 FILLCELL_97_1859 ();
 FILLCELL_X4 FILLCELL_97_1891 ();
 FILLCELL_X2 FILLCELL_97_1895 ();
 FILLCELL_X32 FILLCELL_98_0 ();
 FILLCELL_X32 FILLCELL_98_32 ();
 FILLCELL_X32 FILLCELL_98_64 ();
 FILLCELL_X32 FILLCELL_98_96 ();
 FILLCELL_X32 FILLCELL_98_128 ();
 FILLCELL_X32 FILLCELL_98_160 ();
 FILLCELL_X32 FILLCELL_98_192 ();
 FILLCELL_X32 FILLCELL_98_224 ();
 FILLCELL_X32 FILLCELL_98_256 ();
 FILLCELL_X32 FILLCELL_98_288 ();
 FILLCELL_X4 FILLCELL_98_320 ();
 FILLCELL_X32 FILLCELL_98_327 ();
 FILLCELL_X32 FILLCELL_98_359 ();
 FILLCELL_X32 FILLCELL_98_391 ();
 FILLCELL_X32 FILLCELL_98_423 ();
 FILLCELL_X32 FILLCELL_98_455 ();
 FILLCELL_X32 FILLCELL_98_487 ();
 FILLCELL_X8 FILLCELL_98_519 ();
 FILLCELL_X32 FILLCELL_98_531 ();
 FILLCELL_X32 FILLCELL_98_563 ();
 FILLCELL_X4 FILLCELL_98_595 ();
 FILLCELL_X2 FILLCELL_98_599 ();
 FILLCELL_X1 FILLCELL_98_601 ();
 FILLCELL_X32 FILLCELL_98_604 ();
 FILLCELL_X32 FILLCELL_98_636 ();
 FILLCELL_X32 FILLCELL_98_668 ();
 FILLCELL_X32 FILLCELL_98_700 ();
 FILLCELL_X32 FILLCELL_98_732 ();
 FILLCELL_X32 FILLCELL_98_764 ();
 FILLCELL_X32 FILLCELL_98_796 ();
 FILLCELL_X8 FILLCELL_98_828 ();
 FILLCELL_X2 FILLCELL_98_836 ();
 FILLCELL_X1 FILLCELL_98_838 ();
 FILLCELL_X4 FILLCELL_98_841 ();
 FILLCELL_X1 FILLCELL_98_845 ();
 FILLCELL_X32 FILLCELL_98_849 ();
 FILLCELL_X32 FILLCELL_98_881 ();
 FILLCELL_X32 FILLCELL_98_913 ();
 FILLCELL_X16 FILLCELL_98_945 ();
 FILLCELL_X8 FILLCELL_98_961 ();
 FILLCELL_X4 FILLCELL_98_969 ();
 FILLCELL_X32 FILLCELL_98_976 ();
 FILLCELL_X32 FILLCELL_98_1008 ();
 FILLCELL_X32 FILLCELL_98_1040 ();
 FILLCELL_X32 FILLCELL_98_1072 ();
 FILLCELL_X32 FILLCELL_98_1104 ();
 FILLCELL_X32 FILLCELL_98_1136 ();
 FILLCELL_X32 FILLCELL_98_1168 ();
 FILLCELL_X32 FILLCELL_98_1200 ();
 FILLCELL_X32 FILLCELL_98_1232 ();
 FILLCELL_X32 FILLCELL_98_1264 ();
 FILLCELL_X32 FILLCELL_98_1296 ();
 FILLCELL_X32 FILLCELL_98_1328 ();
 FILLCELL_X32 FILLCELL_98_1360 ();
 FILLCELL_X32 FILLCELL_98_1392 ();
 FILLCELL_X32 FILLCELL_98_1424 ();
 FILLCELL_X32 FILLCELL_98_1456 ();
 FILLCELL_X32 FILLCELL_98_1488 ();
 FILLCELL_X32 FILLCELL_98_1520 ();
 FILLCELL_X32 FILLCELL_98_1552 ();
 FILLCELL_X32 FILLCELL_98_1584 ();
 FILLCELL_X32 FILLCELL_98_1616 ();
 FILLCELL_X32 FILLCELL_98_1648 ();
 FILLCELL_X32 FILLCELL_98_1680 ();
 FILLCELL_X32 FILLCELL_98_1712 ();
 FILLCELL_X32 FILLCELL_98_1744 ();
 FILLCELL_X32 FILLCELL_98_1776 ();
 FILLCELL_X32 FILLCELL_98_1808 ();
 FILLCELL_X32 FILLCELL_98_1840 ();
 FILLCELL_X16 FILLCELL_98_1872 ();
 FILLCELL_X8 FILLCELL_98_1888 ();
 FILLCELL_X1 FILLCELL_98_1896 ();
 FILLCELL_X32 FILLCELL_99_0 ();
 FILLCELL_X32 FILLCELL_99_32 ();
 FILLCELL_X32 FILLCELL_99_64 ();
 FILLCELL_X32 FILLCELL_99_96 ();
 FILLCELL_X32 FILLCELL_99_128 ();
 FILLCELL_X32 FILLCELL_99_160 ();
 FILLCELL_X16 FILLCELL_99_192 ();
 FILLCELL_X4 FILLCELL_99_208 ();
 FILLCELL_X2 FILLCELL_99_212 ();
 FILLCELL_X32 FILLCELL_99_217 ();
 FILLCELL_X32 FILLCELL_99_249 ();
 FILLCELL_X32 FILLCELL_99_281 ();
 FILLCELL_X32 FILLCELL_99_313 ();
 FILLCELL_X32 FILLCELL_99_345 ();
 FILLCELL_X32 FILLCELL_99_377 ();
 FILLCELL_X32 FILLCELL_99_409 ();
 FILLCELL_X32 FILLCELL_99_441 ();
 FILLCELL_X32 FILLCELL_99_473 ();
 FILLCELL_X32 FILLCELL_99_505 ();
 FILLCELL_X16 FILLCELL_99_537 ();
 FILLCELL_X8 FILLCELL_99_553 ();
 FILLCELL_X1 FILLCELL_99_561 ();
 FILLCELL_X32 FILLCELL_99_566 ();
 FILLCELL_X4 FILLCELL_99_598 ();
 FILLCELL_X32 FILLCELL_99_607 ();
 FILLCELL_X32 FILLCELL_99_639 ();
 FILLCELL_X32 FILLCELL_99_671 ();
 FILLCELL_X32 FILLCELL_99_703 ();
 FILLCELL_X32 FILLCELL_99_735 ();
 FILLCELL_X32 FILLCELL_99_767 ();
 FILLCELL_X32 FILLCELL_99_799 ();
 FILLCELL_X32 FILLCELL_99_831 ();
 FILLCELL_X32 FILLCELL_99_863 ();
 FILLCELL_X32 FILLCELL_99_895 ();
 FILLCELL_X32 FILLCELL_99_927 ();
 FILLCELL_X32 FILLCELL_99_959 ();
 FILLCELL_X32 FILLCELL_99_991 ();
 FILLCELL_X32 FILLCELL_99_1023 ();
 FILLCELL_X32 FILLCELL_99_1055 ();
 FILLCELL_X32 FILLCELL_99_1087 ();
 FILLCELL_X32 FILLCELL_99_1119 ();
 FILLCELL_X32 FILLCELL_99_1151 ();
 FILLCELL_X32 FILLCELL_99_1183 ();
 FILLCELL_X32 FILLCELL_99_1215 ();
 FILLCELL_X32 FILLCELL_99_1247 ();
 FILLCELL_X32 FILLCELL_99_1279 ();
 FILLCELL_X32 FILLCELL_99_1311 ();
 FILLCELL_X32 FILLCELL_99_1343 ();
 FILLCELL_X32 FILLCELL_99_1375 ();
 FILLCELL_X32 FILLCELL_99_1407 ();
 FILLCELL_X32 FILLCELL_99_1439 ();
 FILLCELL_X32 FILLCELL_99_1471 ();
 FILLCELL_X32 FILLCELL_99_1503 ();
 FILLCELL_X32 FILLCELL_99_1535 ();
 FILLCELL_X32 FILLCELL_99_1567 ();
 FILLCELL_X32 FILLCELL_99_1599 ();
 FILLCELL_X32 FILLCELL_99_1631 ();
 FILLCELL_X32 FILLCELL_99_1663 ();
 FILLCELL_X32 FILLCELL_99_1695 ();
 FILLCELL_X32 FILLCELL_99_1727 ();
 FILLCELL_X32 FILLCELL_99_1759 ();
 FILLCELL_X32 FILLCELL_99_1791 ();
 FILLCELL_X32 FILLCELL_99_1823 ();
 FILLCELL_X32 FILLCELL_99_1855 ();
 FILLCELL_X8 FILLCELL_99_1887 ();
 FILLCELL_X2 FILLCELL_99_1895 ();
 FILLCELL_X32 FILLCELL_100_0 ();
 FILLCELL_X32 FILLCELL_100_32 ();
 FILLCELL_X32 FILLCELL_100_64 ();
 FILLCELL_X32 FILLCELL_100_96 ();
 FILLCELL_X32 FILLCELL_100_128 ();
 FILLCELL_X32 FILLCELL_100_160 ();
 FILLCELL_X32 FILLCELL_100_192 ();
 FILLCELL_X32 FILLCELL_100_224 ();
 FILLCELL_X32 FILLCELL_100_256 ();
 FILLCELL_X32 FILLCELL_100_288 ();
 FILLCELL_X32 FILLCELL_100_320 ();
 FILLCELL_X16 FILLCELL_100_352 ();
 FILLCELL_X2 FILLCELL_100_368 ();
 FILLCELL_X1 FILLCELL_100_370 ();
 FILLCELL_X32 FILLCELL_100_373 ();
 FILLCELL_X32 FILLCELL_100_405 ();
 FILLCELL_X1 FILLCELL_100_437 ();
 FILLCELL_X32 FILLCELL_100_441 ();
 FILLCELL_X32 FILLCELL_100_473 ();
 FILLCELL_X32 FILLCELL_100_505 ();
 FILLCELL_X32 FILLCELL_100_537 ();
 FILLCELL_X32 FILLCELL_100_569 ();
 FILLCELL_X32 FILLCELL_100_601 ();
 FILLCELL_X32 FILLCELL_100_633 ();
 FILLCELL_X32 FILLCELL_100_665 ();
 FILLCELL_X32 FILLCELL_100_697 ();
 FILLCELL_X32 FILLCELL_100_729 ();
 FILLCELL_X32 FILLCELL_100_761 ();
 FILLCELL_X32 FILLCELL_100_793 ();
 FILLCELL_X32 FILLCELL_100_825 ();
 FILLCELL_X32 FILLCELL_100_857 ();
 FILLCELL_X32 FILLCELL_100_889 ();
 FILLCELL_X32 FILLCELL_100_921 ();
 FILLCELL_X32 FILLCELL_100_953 ();
 FILLCELL_X32 FILLCELL_100_985 ();
 FILLCELL_X32 FILLCELL_100_1017 ();
 FILLCELL_X32 FILLCELL_100_1049 ();
 FILLCELL_X32 FILLCELL_100_1081 ();
 FILLCELL_X32 FILLCELL_100_1113 ();
 FILLCELL_X32 FILLCELL_100_1145 ();
 FILLCELL_X32 FILLCELL_100_1177 ();
 FILLCELL_X32 FILLCELL_100_1209 ();
 FILLCELL_X32 FILLCELL_100_1241 ();
 FILLCELL_X32 FILLCELL_100_1273 ();
 FILLCELL_X32 FILLCELL_100_1305 ();
 FILLCELL_X32 FILLCELL_100_1337 ();
 FILLCELL_X32 FILLCELL_100_1369 ();
 FILLCELL_X32 FILLCELL_100_1401 ();
 FILLCELL_X32 FILLCELL_100_1433 ();
 FILLCELL_X32 FILLCELL_100_1465 ();
 FILLCELL_X32 FILLCELL_100_1497 ();
 FILLCELL_X32 FILLCELL_100_1529 ();
 FILLCELL_X32 FILLCELL_100_1561 ();
 FILLCELL_X32 FILLCELL_100_1593 ();
 FILLCELL_X32 FILLCELL_100_1625 ();
 FILLCELL_X32 FILLCELL_100_1657 ();
 FILLCELL_X32 FILLCELL_100_1689 ();
 FILLCELL_X32 FILLCELL_100_1721 ();
 FILLCELL_X32 FILLCELL_100_1753 ();
 FILLCELL_X32 FILLCELL_100_1785 ();
 FILLCELL_X32 FILLCELL_100_1817 ();
 FILLCELL_X32 FILLCELL_100_1849 ();
 FILLCELL_X16 FILLCELL_100_1881 ();
 FILLCELL_X32 FILLCELL_101_0 ();
 FILLCELL_X32 FILLCELL_101_32 ();
 FILLCELL_X32 FILLCELL_101_64 ();
 FILLCELL_X32 FILLCELL_101_96 ();
 FILLCELL_X32 FILLCELL_101_128 ();
 FILLCELL_X16 FILLCELL_101_160 ();
 FILLCELL_X2 FILLCELL_101_176 ();
 FILLCELL_X32 FILLCELL_101_183 ();
 FILLCELL_X32 FILLCELL_101_215 ();
 FILLCELL_X32 FILLCELL_101_247 ();
 FILLCELL_X32 FILLCELL_101_279 ();
 FILLCELL_X32 FILLCELL_101_311 ();
 FILLCELL_X32 FILLCELL_101_343 ();
 FILLCELL_X32 FILLCELL_101_375 ();
 FILLCELL_X32 FILLCELL_101_407 ();
 FILLCELL_X32 FILLCELL_101_439 ();
 FILLCELL_X32 FILLCELL_101_471 ();
 FILLCELL_X32 FILLCELL_101_503 ();
 FILLCELL_X32 FILLCELL_101_535 ();
 FILLCELL_X32 FILLCELL_101_567 ();
 FILLCELL_X32 FILLCELL_101_599 ();
 FILLCELL_X32 FILLCELL_101_631 ();
 FILLCELL_X32 FILLCELL_101_663 ();
 FILLCELL_X32 FILLCELL_101_695 ();
 FILLCELL_X32 FILLCELL_101_727 ();
 FILLCELL_X32 FILLCELL_101_759 ();
 FILLCELL_X8 FILLCELL_101_791 ();
 FILLCELL_X32 FILLCELL_101_802 ();
 FILLCELL_X32 FILLCELL_101_834 ();
 FILLCELL_X32 FILLCELL_101_866 ();
 FILLCELL_X32 FILLCELL_101_898 ();
 FILLCELL_X32 FILLCELL_101_930 ();
 FILLCELL_X32 FILLCELL_101_962 ();
 FILLCELL_X32 FILLCELL_101_994 ();
 FILLCELL_X32 FILLCELL_101_1026 ();
 FILLCELL_X32 FILLCELL_101_1058 ();
 FILLCELL_X32 FILLCELL_101_1090 ();
 FILLCELL_X32 FILLCELL_101_1122 ();
 FILLCELL_X32 FILLCELL_101_1154 ();
 FILLCELL_X32 FILLCELL_101_1186 ();
 FILLCELL_X32 FILLCELL_101_1218 ();
 FILLCELL_X32 FILLCELL_101_1250 ();
 FILLCELL_X32 FILLCELL_101_1282 ();
 FILLCELL_X32 FILLCELL_101_1314 ();
 FILLCELL_X32 FILLCELL_101_1346 ();
 FILLCELL_X32 FILLCELL_101_1378 ();
 FILLCELL_X32 FILLCELL_101_1410 ();
 FILLCELL_X32 FILLCELL_101_1442 ();
 FILLCELL_X32 FILLCELL_101_1474 ();
 FILLCELL_X32 FILLCELL_101_1506 ();
 FILLCELL_X32 FILLCELL_101_1538 ();
 FILLCELL_X32 FILLCELL_101_1570 ();
 FILLCELL_X32 FILLCELL_101_1602 ();
 FILLCELL_X32 FILLCELL_101_1634 ();
 FILLCELL_X32 FILLCELL_101_1666 ();
 FILLCELL_X32 FILLCELL_101_1698 ();
 FILLCELL_X32 FILLCELL_101_1730 ();
 FILLCELL_X32 FILLCELL_101_1762 ();
 FILLCELL_X32 FILLCELL_101_1794 ();
 FILLCELL_X32 FILLCELL_101_1826 ();
 FILLCELL_X32 FILLCELL_101_1858 ();
 FILLCELL_X4 FILLCELL_101_1890 ();
 FILLCELL_X2 FILLCELL_101_1894 ();
 FILLCELL_X1 FILLCELL_101_1896 ();
 FILLCELL_X32 FILLCELL_102_0 ();
 FILLCELL_X32 FILLCELL_102_32 ();
 FILLCELL_X32 FILLCELL_102_64 ();
 FILLCELL_X32 FILLCELL_102_96 ();
 FILLCELL_X32 FILLCELL_102_128 ();
 FILLCELL_X32 FILLCELL_102_160 ();
 FILLCELL_X32 FILLCELL_102_192 ();
 FILLCELL_X32 FILLCELL_102_224 ();
 FILLCELL_X32 FILLCELL_102_256 ();
 FILLCELL_X16 FILLCELL_102_288 ();
 FILLCELL_X4 FILLCELL_102_304 ();
 FILLCELL_X2 FILLCELL_102_308 ();
 FILLCELL_X1 FILLCELL_102_310 ();
 FILLCELL_X32 FILLCELL_102_314 ();
 FILLCELL_X32 FILLCELL_102_346 ();
 FILLCELL_X32 FILLCELL_102_378 ();
 FILLCELL_X16 FILLCELL_102_410 ();
 FILLCELL_X2 FILLCELL_102_426 ();
 FILLCELL_X32 FILLCELL_102_431 ();
 FILLCELL_X32 FILLCELL_102_463 ();
 FILLCELL_X32 FILLCELL_102_495 ();
 FILLCELL_X32 FILLCELL_102_527 ();
 FILLCELL_X32 FILLCELL_102_559 ();
 FILLCELL_X32 FILLCELL_102_591 ();
 FILLCELL_X32 FILLCELL_102_623 ();
 FILLCELL_X32 FILLCELL_102_655 ();
 FILLCELL_X32 FILLCELL_102_687 ();
 FILLCELL_X32 FILLCELL_102_719 ();
 FILLCELL_X32 FILLCELL_102_751 ();
 FILLCELL_X32 FILLCELL_102_783 ();
 FILLCELL_X32 FILLCELL_102_815 ();
 FILLCELL_X32 FILLCELL_102_847 ();
 FILLCELL_X32 FILLCELL_102_879 ();
 FILLCELL_X16 FILLCELL_102_911 ();
 FILLCELL_X4 FILLCELL_102_927 ();
 FILLCELL_X2 FILLCELL_102_931 ();
 FILLCELL_X1 FILLCELL_102_933 ();
 FILLCELL_X8 FILLCELL_102_937 ();
 FILLCELL_X2 FILLCELL_102_945 ();
 FILLCELL_X1 FILLCELL_102_947 ();
 FILLCELL_X32 FILLCELL_102_951 ();
 FILLCELL_X32 FILLCELL_102_983 ();
 FILLCELL_X32 FILLCELL_102_1015 ();
 FILLCELL_X32 FILLCELL_102_1047 ();
 FILLCELL_X32 FILLCELL_102_1079 ();
 FILLCELL_X32 FILLCELL_102_1111 ();
 FILLCELL_X32 FILLCELL_102_1143 ();
 FILLCELL_X32 FILLCELL_102_1175 ();
 FILLCELL_X32 FILLCELL_102_1207 ();
 FILLCELL_X32 FILLCELL_102_1239 ();
 FILLCELL_X32 FILLCELL_102_1271 ();
 FILLCELL_X32 FILLCELL_102_1303 ();
 FILLCELL_X32 FILLCELL_102_1335 ();
 FILLCELL_X32 FILLCELL_102_1367 ();
 FILLCELL_X32 FILLCELL_102_1399 ();
 FILLCELL_X32 FILLCELL_102_1431 ();
 FILLCELL_X32 FILLCELL_102_1463 ();
 FILLCELL_X32 FILLCELL_102_1495 ();
 FILLCELL_X32 FILLCELL_102_1527 ();
 FILLCELL_X32 FILLCELL_102_1559 ();
 FILLCELL_X32 FILLCELL_102_1591 ();
 FILLCELL_X32 FILLCELL_102_1623 ();
 FILLCELL_X32 FILLCELL_102_1655 ();
 FILLCELL_X32 FILLCELL_102_1687 ();
 FILLCELL_X32 FILLCELL_102_1719 ();
 FILLCELL_X32 FILLCELL_102_1751 ();
 FILLCELL_X32 FILLCELL_102_1783 ();
 FILLCELL_X32 FILLCELL_102_1815 ();
 FILLCELL_X32 FILLCELL_102_1847 ();
 FILLCELL_X16 FILLCELL_102_1879 ();
 FILLCELL_X2 FILLCELL_102_1895 ();
 FILLCELL_X32 FILLCELL_103_0 ();
 FILLCELL_X16 FILLCELL_103_32 ();
 FILLCELL_X4 FILLCELL_103_48 ();
 FILLCELL_X1 FILLCELL_103_52 ();
 FILLCELL_X32 FILLCELL_103_70 ();
 FILLCELL_X32 FILLCELL_103_102 ();
 FILLCELL_X32 FILLCELL_103_137 ();
 FILLCELL_X32 FILLCELL_103_169 ();
 FILLCELL_X32 FILLCELL_103_201 ();
 FILLCELL_X32 FILLCELL_103_233 ();
 FILLCELL_X32 FILLCELL_103_265 ();
 FILLCELL_X32 FILLCELL_103_297 ();
 FILLCELL_X32 FILLCELL_103_329 ();
 FILLCELL_X32 FILLCELL_103_361 ();
 FILLCELL_X32 FILLCELL_103_393 ();
 FILLCELL_X32 FILLCELL_103_425 ();
 FILLCELL_X4 FILLCELL_103_457 ();
 FILLCELL_X2 FILLCELL_103_461 ();
 FILLCELL_X1 FILLCELL_103_463 ();
 FILLCELL_X16 FILLCELL_103_466 ();
 FILLCELL_X8 FILLCELL_103_482 ();
 FILLCELL_X4 FILLCELL_103_490 ();
 FILLCELL_X32 FILLCELL_103_499 ();
 FILLCELL_X32 FILLCELL_103_531 ();
 FILLCELL_X32 FILLCELL_103_563 ();
 FILLCELL_X32 FILLCELL_103_595 ();
 FILLCELL_X32 FILLCELL_103_627 ();
 FILLCELL_X32 FILLCELL_103_659 ();
 FILLCELL_X32 FILLCELL_103_691 ();
 FILLCELL_X4 FILLCELL_103_723 ();
 FILLCELL_X1 FILLCELL_103_727 ();
 FILLCELL_X32 FILLCELL_103_735 ();
 FILLCELL_X32 FILLCELL_103_767 ();
 FILLCELL_X32 FILLCELL_103_799 ();
 FILLCELL_X32 FILLCELL_103_831 ();
 FILLCELL_X32 FILLCELL_103_863 ();
 FILLCELL_X32 FILLCELL_103_895 ();
 FILLCELL_X16 FILLCELL_103_927 ();
 FILLCELL_X32 FILLCELL_103_948 ();
 FILLCELL_X32 FILLCELL_103_980 ();
 FILLCELL_X32 FILLCELL_103_1012 ();
 FILLCELL_X32 FILLCELL_103_1044 ();
 FILLCELL_X32 FILLCELL_103_1076 ();
 FILLCELL_X32 FILLCELL_103_1108 ();
 FILLCELL_X32 FILLCELL_103_1140 ();
 FILLCELL_X32 FILLCELL_103_1172 ();
 FILLCELL_X32 FILLCELL_103_1204 ();
 FILLCELL_X32 FILLCELL_103_1236 ();
 FILLCELL_X32 FILLCELL_103_1268 ();
 FILLCELL_X32 FILLCELL_103_1300 ();
 FILLCELL_X32 FILLCELL_103_1332 ();
 FILLCELL_X32 FILLCELL_103_1364 ();
 FILLCELL_X32 FILLCELL_103_1396 ();
 FILLCELL_X32 FILLCELL_103_1428 ();
 FILLCELL_X32 FILLCELL_103_1460 ();
 FILLCELL_X32 FILLCELL_103_1492 ();
 FILLCELL_X32 FILLCELL_103_1524 ();
 FILLCELL_X32 FILLCELL_103_1556 ();
 FILLCELL_X32 FILLCELL_103_1588 ();
 FILLCELL_X32 FILLCELL_103_1620 ();
 FILLCELL_X32 FILLCELL_103_1652 ();
 FILLCELL_X32 FILLCELL_103_1684 ();
 FILLCELL_X32 FILLCELL_103_1716 ();
 FILLCELL_X32 FILLCELL_103_1748 ();
 FILLCELL_X32 FILLCELL_103_1780 ();
 FILLCELL_X32 FILLCELL_103_1812 ();
 FILLCELL_X32 FILLCELL_103_1844 ();
 FILLCELL_X16 FILLCELL_103_1876 ();
 FILLCELL_X4 FILLCELL_103_1892 ();
 FILLCELL_X1 FILLCELL_103_1896 ();
 FILLCELL_X32 FILLCELL_104_0 ();
 FILLCELL_X32 FILLCELL_104_32 ();
 FILLCELL_X32 FILLCELL_104_64 ();
 FILLCELL_X32 FILLCELL_104_96 ();
 FILLCELL_X2 FILLCELL_104_128 ();
 FILLCELL_X1 FILLCELL_104_130 ();
 FILLCELL_X32 FILLCELL_104_135 ();
 FILLCELL_X32 FILLCELL_104_167 ();
 FILLCELL_X32 FILLCELL_104_199 ();
 FILLCELL_X32 FILLCELL_104_231 ();
 FILLCELL_X32 FILLCELL_104_263 ();
 FILLCELL_X32 FILLCELL_104_295 ();
 FILLCELL_X32 FILLCELL_104_327 ();
 FILLCELL_X32 FILLCELL_104_359 ();
 FILLCELL_X32 FILLCELL_104_391 ();
 FILLCELL_X16 FILLCELL_104_423 ();
 FILLCELL_X8 FILLCELL_104_439 ();
 FILLCELL_X2 FILLCELL_104_447 ();
 FILLCELL_X16 FILLCELL_104_453 ();
 FILLCELL_X1 FILLCELL_104_469 ();
 FILLCELL_X32 FILLCELL_104_473 ();
 FILLCELL_X32 FILLCELL_104_505 ();
 FILLCELL_X32 FILLCELL_104_537 ();
 FILLCELL_X16 FILLCELL_104_569 ();
 FILLCELL_X8 FILLCELL_104_585 ();
 FILLCELL_X4 FILLCELL_104_593 ();
 FILLCELL_X1 FILLCELL_104_597 ();
 FILLCELL_X32 FILLCELL_104_601 ();
 FILLCELL_X32 FILLCELL_104_633 ();
 FILLCELL_X32 FILLCELL_104_665 ();
 FILLCELL_X32 FILLCELL_104_697 ();
 FILLCELL_X32 FILLCELL_104_729 ();
 FILLCELL_X32 FILLCELL_104_761 ();
 FILLCELL_X32 FILLCELL_104_793 ();
 FILLCELL_X16 FILLCELL_104_825 ();
 FILLCELL_X8 FILLCELL_104_841 ();
 FILLCELL_X1 FILLCELL_104_849 ();
 FILLCELL_X32 FILLCELL_104_858 ();
 FILLCELL_X32 FILLCELL_104_890 ();
 FILLCELL_X32 FILLCELL_104_922 ();
 FILLCELL_X32 FILLCELL_104_954 ();
 FILLCELL_X32 FILLCELL_104_986 ();
 FILLCELL_X32 FILLCELL_104_1018 ();
 FILLCELL_X32 FILLCELL_104_1050 ();
 FILLCELL_X32 FILLCELL_104_1082 ();
 FILLCELL_X32 FILLCELL_104_1114 ();
 FILLCELL_X32 FILLCELL_104_1146 ();
 FILLCELL_X32 FILLCELL_104_1178 ();
 FILLCELL_X32 FILLCELL_104_1210 ();
 FILLCELL_X32 FILLCELL_104_1242 ();
 FILLCELL_X32 FILLCELL_104_1274 ();
 FILLCELL_X32 FILLCELL_104_1306 ();
 FILLCELL_X32 FILLCELL_104_1338 ();
 FILLCELL_X32 FILLCELL_104_1370 ();
 FILLCELL_X32 FILLCELL_104_1402 ();
 FILLCELL_X32 FILLCELL_104_1434 ();
 FILLCELL_X32 FILLCELL_104_1466 ();
 FILLCELL_X32 FILLCELL_104_1498 ();
 FILLCELL_X32 FILLCELL_104_1530 ();
 FILLCELL_X32 FILLCELL_104_1562 ();
 FILLCELL_X32 FILLCELL_104_1594 ();
 FILLCELL_X32 FILLCELL_104_1626 ();
 FILLCELL_X32 FILLCELL_104_1658 ();
 FILLCELL_X32 FILLCELL_104_1690 ();
 FILLCELL_X32 FILLCELL_104_1722 ();
 FILLCELL_X32 FILLCELL_104_1754 ();
 FILLCELL_X32 FILLCELL_104_1786 ();
 FILLCELL_X32 FILLCELL_104_1818 ();
 FILLCELL_X32 FILLCELL_104_1850 ();
 FILLCELL_X8 FILLCELL_104_1882 ();
 FILLCELL_X4 FILLCELL_104_1890 ();
 FILLCELL_X2 FILLCELL_104_1894 ();
 FILLCELL_X1 FILLCELL_104_1896 ();
 FILLCELL_X32 FILLCELL_105_0 ();
 FILLCELL_X32 FILLCELL_105_32 ();
 FILLCELL_X32 FILLCELL_105_64 ();
 FILLCELL_X32 FILLCELL_105_96 ();
 FILLCELL_X4 FILLCELL_105_128 ();
 FILLCELL_X1 FILLCELL_105_132 ();
 FILLCELL_X16 FILLCELL_105_137 ();
 FILLCELL_X4 FILLCELL_105_153 ();
 FILLCELL_X1 FILLCELL_105_157 ();
 FILLCELL_X32 FILLCELL_105_165 ();
 FILLCELL_X32 FILLCELL_105_197 ();
 FILLCELL_X32 FILLCELL_105_229 ();
 FILLCELL_X32 FILLCELL_105_261 ();
 FILLCELL_X4 FILLCELL_105_293 ();
 FILLCELL_X2 FILLCELL_105_297 ();
 FILLCELL_X32 FILLCELL_105_303 ();
 FILLCELL_X32 FILLCELL_105_335 ();
 FILLCELL_X8 FILLCELL_105_367 ();
 FILLCELL_X4 FILLCELL_105_375 ();
 FILLCELL_X1 FILLCELL_105_379 ();
 FILLCELL_X32 FILLCELL_105_383 ();
 FILLCELL_X32 FILLCELL_105_415 ();
 FILLCELL_X32 FILLCELL_105_447 ();
 FILLCELL_X32 FILLCELL_105_479 ();
 FILLCELL_X32 FILLCELL_105_511 ();
 FILLCELL_X32 FILLCELL_105_543 ();
 FILLCELL_X32 FILLCELL_105_575 ();
 FILLCELL_X32 FILLCELL_105_607 ();
 FILLCELL_X32 FILLCELL_105_639 ();
 FILLCELL_X32 FILLCELL_105_671 ();
 FILLCELL_X16 FILLCELL_105_703 ();
 FILLCELL_X32 FILLCELL_105_736 ();
 FILLCELL_X32 FILLCELL_105_768 ();
 FILLCELL_X32 FILLCELL_105_800 ();
 FILLCELL_X2 FILLCELL_105_832 ();
 FILLCELL_X32 FILLCELL_105_837 ();
 FILLCELL_X32 FILLCELL_105_869 ();
 FILLCELL_X16 FILLCELL_105_901 ();
 FILLCELL_X2 FILLCELL_105_917 ();
 FILLCELL_X32 FILLCELL_105_923 ();
 FILLCELL_X32 FILLCELL_105_955 ();
 FILLCELL_X32 FILLCELL_105_987 ();
 FILLCELL_X32 FILLCELL_105_1019 ();
 FILLCELL_X32 FILLCELL_105_1051 ();
 FILLCELL_X16 FILLCELL_105_1083 ();
 FILLCELL_X2 FILLCELL_105_1099 ();
 FILLCELL_X32 FILLCELL_105_1108 ();
 FILLCELL_X32 FILLCELL_105_1140 ();
 FILLCELL_X32 FILLCELL_105_1172 ();
 FILLCELL_X32 FILLCELL_105_1204 ();
 FILLCELL_X32 FILLCELL_105_1236 ();
 FILLCELL_X32 FILLCELL_105_1268 ();
 FILLCELL_X32 FILLCELL_105_1300 ();
 FILLCELL_X32 FILLCELL_105_1332 ();
 FILLCELL_X32 FILLCELL_105_1364 ();
 FILLCELL_X32 FILLCELL_105_1396 ();
 FILLCELL_X32 FILLCELL_105_1428 ();
 FILLCELL_X32 FILLCELL_105_1460 ();
 FILLCELL_X32 FILLCELL_105_1492 ();
 FILLCELL_X32 FILLCELL_105_1524 ();
 FILLCELL_X32 FILLCELL_105_1556 ();
 FILLCELL_X32 FILLCELL_105_1588 ();
 FILLCELL_X32 FILLCELL_105_1620 ();
 FILLCELL_X32 FILLCELL_105_1652 ();
 FILLCELL_X32 FILLCELL_105_1684 ();
 FILLCELL_X32 FILLCELL_105_1716 ();
 FILLCELL_X32 FILLCELL_105_1748 ();
 FILLCELL_X32 FILLCELL_105_1780 ();
 FILLCELL_X32 FILLCELL_105_1812 ();
 FILLCELL_X32 FILLCELL_105_1844 ();
 FILLCELL_X16 FILLCELL_105_1876 ();
 FILLCELL_X4 FILLCELL_105_1892 ();
 FILLCELL_X1 FILLCELL_105_1896 ();
 FILLCELL_X32 FILLCELL_106_0 ();
 FILLCELL_X32 FILLCELL_106_32 ();
 FILLCELL_X32 FILLCELL_106_64 ();
 FILLCELL_X32 FILLCELL_106_96 ();
 FILLCELL_X32 FILLCELL_106_128 ();
 FILLCELL_X32 FILLCELL_106_160 ();
 FILLCELL_X32 FILLCELL_106_192 ();
 FILLCELL_X32 FILLCELL_106_224 ();
 FILLCELL_X32 FILLCELL_106_256 ();
 FILLCELL_X8 FILLCELL_106_288 ();
 FILLCELL_X2 FILLCELL_106_296 ();
 FILLCELL_X32 FILLCELL_106_302 ();
 FILLCELL_X32 FILLCELL_106_334 ();
 FILLCELL_X4 FILLCELL_106_366 ();
 FILLCELL_X16 FILLCELL_106_375 ();
 FILLCELL_X8 FILLCELL_106_391 ();
 FILLCELL_X4 FILLCELL_106_399 ();
 FILLCELL_X32 FILLCELL_106_406 ();
 FILLCELL_X32 FILLCELL_106_438 ();
 FILLCELL_X32 FILLCELL_106_470 ();
 FILLCELL_X32 FILLCELL_106_502 ();
 FILLCELL_X32 FILLCELL_106_534 ();
 FILLCELL_X32 FILLCELL_106_566 ();
 FILLCELL_X32 FILLCELL_106_598 ();
 FILLCELL_X32 FILLCELL_106_630 ();
 FILLCELL_X32 FILLCELL_106_662 ();
 FILLCELL_X32 FILLCELL_106_694 ();
 FILLCELL_X32 FILLCELL_106_726 ();
 FILLCELL_X32 FILLCELL_106_758 ();
 FILLCELL_X32 FILLCELL_106_790 ();
 FILLCELL_X32 FILLCELL_106_822 ();
 FILLCELL_X32 FILLCELL_106_854 ();
 FILLCELL_X32 FILLCELL_106_886 ();
 FILLCELL_X32 FILLCELL_106_918 ();
 FILLCELL_X32 FILLCELL_106_950 ();
 FILLCELL_X32 FILLCELL_106_982 ();
 FILLCELL_X32 FILLCELL_106_1014 ();
 FILLCELL_X8 FILLCELL_106_1046 ();
 FILLCELL_X1 FILLCELL_106_1054 ();
 FILLCELL_X32 FILLCELL_106_1058 ();
 FILLCELL_X16 FILLCELL_106_1090 ();
 FILLCELL_X8 FILLCELL_106_1106 ();
 FILLCELL_X1 FILLCELL_106_1114 ();
 FILLCELL_X32 FILLCELL_106_1120 ();
 FILLCELL_X32 FILLCELL_106_1152 ();
 FILLCELL_X32 FILLCELL_106_1184 ();
 FILLCELL_X32 FILLCELL_106_1216 ();
 FILLCELL_X32 FILLCELL_106_1248 ();
 FILLCELL_X32 FILLCELL_106_1280 ();
 FILLCELL_X32 FILLCELL_106_1312 ();
 FILLCELL_X32 FILLCELL_106_1344 ();
 FILLCELL_X32 FILLCELL_106_1376 ();
 FILLCELL_X32 FILLCELL_106_1408 ();
 FILLCELL_X32 FILLCELL_106_1440 ();
 FILLCELL_X32 FILLCELL_106_1472 ();
 FILLCELL_X32 FILLCELL_106_1504 ();
 FILLCELL_X32 FILLCELL_106_1536 ();
 FILLCELL_X32 FILLCELL_106_1568 ();
 FILLCELL_X32 FILLCELL_106_1600 ();
 FILLCELL_X32 FILLCELL_106_1632 ();
 FILLCELL_X32 FILLCELL_106_1664 ();
 FILLCELL_X32 FILLCELL_106_1696 ();
 FILLCELL_X32 FILLCELL_106_1728 ();
 FILLCELL_X32 FILLCELL_106_1760 ();
 FILLCELL_X32 FILLCELL_106_1792 ();
 FILLCELL_X32 FILLCELL_106_1824 ();
 FILLCELL_X32 FILLCELL_106_1856 ();
 FILLCELL_X8 FILLCELL_106_1888 ();
 FILLCELL_X1 FILLCELL_106_1896 ();
 FILLCELL_X32 FILLCELL_107_0 ();
 FILLCELL_X32 FILLCELL_107_32 ();
 FILLCELL_X32 FILLCELL_107_64 ();
 FILLCELL_X32 FILLCELL_107_96 ();
 FILLCELL_X32 FILLCELL_107_128 ();
 FILLCELL_X32 FILLCELL_107_160 ();
 FILLCELL_X32 FILLCELL_107_192 ();
 FILLCELL_X32 FILLCELL_107_224 ();
 FILLCELL_X32 FILLCELL_107_256 ();
 FILLCELL_X32 FILLCELL_107_288 ();
 FILLCELL_X32 FILLCELL_107_320 ();
 FILLCELL_X32 FILLCELL_107_352 ();
 FILLCELL_X32 FILLCELL_107_384 ();
 FILLCELL_X32 FILLCELL_107_416 ();
 FILLCELL_X32 FILLCELL_107_448 ();
 FILLCELL_X32 FILLCELL_107_480 ();
 FILLCELL_X32 FILLCELL_107_512 ();
 FILLCELL_X32 FILLCELL_107_544 ();
 FILLCELL_X32 FILLCELL_107_576 ();
 FILLCELL_X32 FILLCELL_107_608 ();
 FILLCELL_X32 FILLCELL_107_640 ();
 FILLCELL_X32 FILLCELL_107_672 ();
 FILLCELL_X32 FILLCELL_107_704 ();
 FILLCELL_X32 FILLCELL_107_736 ();
 FILLCELL_X32 FILLCELL_107_768 ();
 FILLCELL_X32 FILLCELL_107_800 ();
 FILLCELL_X32 FILLCELL_107_832 ();
 FILLCELL_X32 FILLCELL_107_864 ();
 FILLCELL_X32 FILLCELL_107_896 ();
 FILLCELL_X32 FILLCELL_107_928 ();
 FILLCELL_X8 FILLCELL_107_960 ();
 FILLCELL_X2 FILLCELL_107_968 ();
 FILLCELL_X32 FILLCELL_107_972 ();
 FILLCELL_X32 FILLCELL_107_1004 ();
 FILLCELL_X32 FILLCELL_107_1036 ();
 FILLCELL_X32 FILLCELL_107_1068 ();
 FILLCELL_X32 FILLCELL_107_1100 ();
 FILLCELL_X32 FILLCELL_107_1132 ();
 FILLCELL_X32 FILLCELL_107_1164 ();
 FILLCELL_X32 FILLCELL_107_1196 ();
 FILLCELL_X32 FILLCELL_107_1228 ();
 FILLCELL_X32 FILLCELL_107_1260 ();
 FILLCELL_X32 FILLCELL_107_1292 ();
 FILLCELL_X32 FILLCELL_107_1324 ();
 FILLCELL_X32 FILLCELL_107_1356 ();
 FILLCELL_X32 FILLCELL_107_1388 ();
 FILLCELL_X32 FILLCELL_107_1420 ();
 FILLCELL_X32 FILLCELL_107_1452 ();
 FILLCELL_X32 FILLCELL_107_1484 ();
 FILLCELL_X32 FILLCELL_107_1516 ();
 FILLCELL_X32 FILLCELL_107_1548 ();
 FILLCELL_X32 FILLCELL_107_1580 ();
 FILLCELL_X32 FILLCELL_107_1612 ();
 FILLCELL_X32 FILLCELL_107_1644 ();
 FILLCELL_X32 FILLCELL_107_1676 ();
 FILLCELL_X32 FILLCELL_107_1708 ();
 FILLCELL_X32 FILLCELL_107_1740 ();
 FILLCELL_X32 FILLCELL_107_1772 ();
 FILLCELL_X32 FILLCELL_107_1804 ();
 FILLCELL_X32 FILLCELL_107_1836 ();
 FILLCELL_X16 FILLCELL_107_1868 ();
 FILLCELL_X8 FILLCELL_107_1884 ();
 FILLCELL_X4 FILLCELL_107_1892 ();
 FILLCELL_X1 FILLCELL_107_1896 ();
 FILLCELL_X32 FILLCELL_108_0 ();
 FILLCELL_X32 FILLCELL_108_32 ();
 FILLCELL_X32 FILLCELL_108_64 ();
 FILLCELL_X32 FILLCELL_108_96 ();
 FILLCELL_X32 FILLCELL_108_128 ();
 FILLCELL_X32 FILLCELL_108_160 ();
 FILLCELL_X32 FILLCELL_108_192 ();
 FILLCELL_X16 FILLCELL_108_224 ();
 FILLCELL_X8 FILLCELL_108_240 ();
 FILLCELL_X4 FILLCELL_108_248 ();
 FILLCELL_X32 FILLCELL_108_255 ();
 FILLCELL_X32 FILLCELL_108_287 ();
 FILLCELL_X32 FILLCELL_108_319 ();
 FILLCELL_X32 FILLCELL_108_351 ();
 FILLCELL_X32 FILLCELL_108_383 ();
 FILLCELL_X32 FILLCELL_108_415 ();
 FILLCELL_X32 FILLCELL_108_447 ();
 FILLCELL_X32 FILLCELL_108_479 ();
 FILLCELL_X32 FILLCELL_108_511 ();
 FILLCELL_X32 FILLCELL_108_543 ();
 FILLCELL_X32 FILLCELL_108_575 ();
 FILLCELL_X32 FILLCELL_108_607 ();
 FILLCELL_X32 FILLCELL_108_639 ();
 FILLCELL_X32 FILLCELL_108_671 ();
 FILLCELL_X32 FILLCELL_108_703 ();
 FILLCELL_X32 FILLCELL_108_735 ();
 FILLCELL_X32 FILLCELL_108_767 ();
 FILLCELL_X32 FILLCELL_108_799 ();
 FILLCELL_X32 FILLCELL_108_831 ();
 FILLCELL_X32 FILLCELL_108_863 ();
 FILLCELL_X32 FILLCELL_108_895 ();
 FILLCELL_X32 FILLCELL_108_927 ();
 FILLCELL_X32 FILLCELL_108_959 ();
 FILLCELL_X32 FILLCELL_108_991 ();
 FILLCELL_X32 FILLCELL_108_1023 ();
 FILLCELL_X32 FILLCELL_108_1055 ();
 FILLCELL_X32 FILLCELL_108_1087 ();
 FILLCELL_X32 FILLCELL_108_1119 ();
 FILLCELL_X32 FILLCELL_108_1151 ();
 FILLCELL_X32 FILLCELL_108_1183 ();
 FILLCELL_X32 FILLCELL_108_1215 ();
 FILLCELL_X32 FILLCELL_108_1247 ();
 FILLCELL_X32 FILLCELL_108_1279 ();
 FILLCELL_X32 FILLCELL_108_1311 ();
 FILLCELL_X32 FILLCELL_108_1343 ();
 FILLCELL_X32 FILLCELL_108_1375 ();
 FILLCELL_X32 FILLCELL_108_1407 ();
 FILLCELL_X32 FILLCELL_108_1439 ();
 FILLCELL_X32 FILLCELL_108_1471 ();
 FILLCELL_X32 FILLCELL_108_1503 ();
 FILLCELL_X32 FILLCELL_108_1535 ();
 FILLCELL_X32 FILLCELL_108_1567 ();
 FILLCELL_X32 FILLCELL_108_1599 ();
 FILLCELL_X32 FILLCELL_108_1631 ();
 FILLCELL_X32 FILLCELL_108_1663 ();
 FILLCELL_X32 FILLCELL_108_1695 ();
 FILLCELL_X32 FILLCELL_108_1727 ();
 FILLCELL_X32 FILLCELL_108_1759 ();
 FILLCELL_X32 FILLCELL_108_1791 ();
 FILLCELL_X32 FILLCELL_108_1823 ();
 FILLCELL_X32 FILLCELL_108_1855 ();
 FILLCELL_X8 FILLCELL_108_1887 ();
 FILLCELL_X2 FILLCELL_108_1895 ();
 FILLCELL_X32 FILLCELL_109_0 ();
 FILLCELL_X32 FILLCELL_109_32 ();
 FILLCELL_X32 FILLCELL_109_64 ();
 FILLCELL_X32 FILLCELL_109_96 ();
 FILLCELL_X32 FILLCELL_109_128 ();
 FILLCELL_X32 FILLCELL_109_160 ();
 FILLCELL_X32 FILLCELL_109_192 ();
 FILLCELL_X16 FILLCELL_109_224 ();
 FILLCELL_X8 FILLCELL_109_240 ();
 FILLCELL_X2 FILLCELL_109_248 ();
 FILLCELL_X16 FILLCELL_109_261 ();
 FILLCELL_X4 FILLCELL_109_277 ();
 FILLCELL_X2 FILLCELL_109_281 ();
 FILLCELL_X32 FILLCELL_109_286 ();
 FILLCELL_X32 FILLCELL_109_318 ();
 FILLCELL_X2 FILLCELL_109_350 ();
 FILLCELL_X1 FILLCELL_109_352 ();
 FILLCELL_X32 FILLCELL_109_356 ();
 FILLCELL_X32 FILLCELL_109_388 ();
 FILLCELL_X8 FILLCELL_109_420 ();
 FILLCELL_X4 FILLCELL_109_428 ();
 FILLCELL_X2 FILLCELL_109_432 ();
 FILLCELL_X1 FILLCELL_109_434 ();
 FILLCELL_X32 FILLCELL_109_438 ();
 FILLCELL_X32 FILLCELL_109_470 ();
 FILLCELL_X32 FILLCELL_109_502 ();
 FILLCELL_X32 FILLCELL_109_534 ();
 FILLCELL_X32 FILLCELL_109_566 ();
 FILLCELL_X32 FILLCELL_109_598 ();
 FILLCELL_X16 FILLCELL_109_630 ();
 FILLCELL_X2 FILLCELL_109_646 ();
 FILLCELL_X32 FILLCELL_109_652 ();
 FILLCELL_X16 FILLCELL_109_684 ();
 FILLCELL_X2 FILLCELL_109_700 ();
 FILLCELL_X32 FILLCELL_109_704 ();
 FILLCELL_X32 FILLCELL_109_736 ();
 FILLCELL_X32 FILLCELL_109_768 ();
 FILLCELL_X16 FILLCELL_109_800 ();
 FILLCELL_X4 FILLCELL_109_816 ();
 FILLCELL_X2 FILLCELL_109_820 ();
 FILLCELL_X32 FILLCELL_109_826 ();
 FILLCELL_X32 FILLCELL_109_858 ();
 FILLCELL_X32 FILLCELL_109_890 ();
 FILLCELL_X32 FILLCELL_109_922 ();
 FILLCELL_X32 FILLCELL_109_954 ();
 FILLCELL_X32 FILLCELL_109_986 ();
 FILLCELL_X32 FILLCELL_109_1018 ();
 FILLCELL_X32 FILLCELL_109_1050 ();
 FILLCELL_X32 FILLCELL_109_1082 ();
 FILLCELL_X32 FILLCELL_109_1114 ();
 FILLCELL_X32 FILLCELL_109_1146 ();
 FILLCELL_X32 FILLCELL_109_1178 ();
 FILLCELL_X32 FILLCELL_109_1210 ();
 FILLCELL_X32 FILLCELL_109_1242 ();
 FILLCELL_X32 FILLCELL_109_1274 ();
 FILLCELL_X32 FILLCELL_109_1306 ();
 FILLCELL_X32 FILLCELL_109_1338 ();
 FILLCELL_X32 FILLCELL_109_1370 ();
 FILLCELL_X32 FILLCELL_109_1402 ();
 FILLCELL_X32 FILLCELL_109_1434 ();
 FILLCELL_X32 FILLCELL_109_1466 ();
 FILLCELL_X32 FILLCELL_109_1498 ();
 FILLCELL_X32 FILLCELL_109_1530 ();
 FILLCELL_X32 FILLCELL_109_1562 ();
 FILLCELL_X32 FILLCELL_109_1594 ();
 FILLCELL_X32 FILLCELL_109_1626 ();
 FILLCELL_X32 FILLCELL_109_1658 ();
 FILLCELL_X32 FILLCELL_109_1690 ();
 FILLCELL_X32 FILLCELL_109_1722 ();
 FILLCELL_X32 FILLCELL_109_1754 ();
 FILLCELL_X32 FILLCELL_109_1786 ();
 FILLCELL_X32 FILLCELL_109_1818 ();
 FILLCELL_X32 FILLCELL_109_1850 ();
 FILLCELL_X8 FILLCELL_109_1882 ();
 FILLCELL_X4 FILLCELL_109_1890 ();
 FILLCELL_X2 FILLCELL_109_1894 ();
 FILLCELL_X1 FILLCELL_109_1896 ();
 FILLCELL_X32 FILLCELL_110_0 ();
 FILLCELL_X32 FILLCELL_110_32 ();
 FILLCELL_X32 FILLCELL_110_64 ();
 FILLCELL_X32 FILLCELL_110_96 ();
 FILLCELL_X32 FILLCELL_110_128 ();
 FILLCELL_X32 FILLCELL_110_160 ();
 FILLCELL_X32 FILLCELL_110_192 ();
 FILLCELL_X32 FILLCELL_110_224 ();
 FILLCELL_X32 FILLCELL_110_256 ();
 FILLCELL_X16 FILLCELL_110_288 ();
 FILLCELL_X8 FILLCELL_110_304 ();
 FILLCELL_X4 FILLCELL_110_312 ();
 FILLCELL_X32 FILLCELL_110_320 ();
 FILLCELL_X32 FILLCELL_110_352 ();
 FILLCELL_X32 FILLCELL_110_384 ();
 FILLCELL_X32 FILLCELL_110_416 ();
 FILLCELL_X32 FILLCELL_110_448 ();
 FILLCELL_X32 FILLCELL_110_480 ();
 FILLCELL_X16 FILLCELL_110_512 ();
 FILLCELL_X8 FILLCELL_110_528 ();
 FILLCELL_X4 FILLCELL_110_536 ();
 FILLCELL_X1 FILLCELL_110_540 ();
 FILLCELL_X32 FILLCELL_110_544 ();
 FILLCELL_X32 FILLCELL_110_576 ();
 FILLCELL_X32 FILLCELL_110_608 ();
 FILLCELL_X32 FILLCELL_110_640 ();
 FILLCELL_X32 FILLCELL_110_672 ();
 FILLCELL_X32 FILLCELL_110_704 ();
 FILLCELL_X32 FILLCELL_110_736 ();
 FILLCELL_X32 FILLCELL_110_768 ();
 FILLCELL_X32 FILLCELL_110_800 ();
 FILLCELL_X32 FILLCELL_110_832 ();
 FILLCELL_X32 FILLCELL_110_864 ();
 FILLCELL_X32 FILLCELL_110_896 ();
 FILLCELL_X32 FILLCELL_110_928 ();
 FILLCELL_X32 FILLCELL_110_960 ();
 FILLCELL_X8 FILLCELL_110_992 ();
 FILLCELL_X4 FILLCELL_110_1000 ();
 FILLCELL_X32 FILLCELL_110_1010 ();
 FILLCELL_X32 FILLCELL_110_1042 ();
 FILLCELL_X32 FILLCELL_110_1074 ();
 FILLCELL_X32 FILLCELL_110_1106 ();
 FILLCELL_X2 FILLCELL_110_1138 ();
 FILLCELL_X32 FILLCELL_110_1147 ();
 FILLCELL_X32 FILLCELL_110_1179 ();
 FILLCELL_X32 FILLCELL_110_1211 ();
 FILLCELL_X32 FILLCELL_110_1243 ();
 FILLCELL_X32 FILLCELL_110_1275 ();
 FILLCELL_X32 FILLCELL_110_1307 ();
 FILLCELL_X32 FILLCELL_110_1339 ();
 FILLCELL_X32 FILLCELL_110_1371 ();
 FILLCELL_X32 FILLCELL_110_1403 ();
 FILLCELL_X32 FILLCELL_110_1435 ();
 FILLCELL_X32 FILLCELL_110_1467 ();
 FILLCELL_X32 FILLCELL_110_1499 ();
 FILLCELL_X32 FILLCELL_110_1531 ();
 FILLCELL_X32 FILLCELL_110_1563 ();
 FILLCELL_X32 FILLCELL_110_1595 ();
 FILLCELL_X32 FILLCELL_110_1627 ();
 FILLCELL_X32 FILLCELL_110_1659 ();
 FILLCELL_X32 FILLCELL_110_1691 ();
 FILLCELL_X32 FILLCELL_110_1723 ();
 FILLCELL_X32 FILLCELL_110_1755 ();
 FILLCELL_X32 FILLCELL_110_1787 ();
 FILLCELL_X32 FILLCELL_110_1819 ();
 FILLCELL_X32 FILLCELL_110_1851 ();
 FILLCELL_X8 FILLCELL_110_1883 ();
 FILLCELL_X4 FILLCELL_110_1891 ();
 FILLCELL_X2 FILLCELL_110_1895 ();
 FILLCELL_X32 FILLCELL_111_0 ();
 FILLCELL_X32 FILLCELL_111_32 ();
 FILLCELL_X32 FILLCELL_111_64 ();
 FILLCELL_X32 FILLCELL_111_96 ();
 FILLCELL_X32 FILLCELL_111_128 ();
 FILLCELL_X32 FILLCELL_111_160 ();
 FILLCELL_X32 FILLCELL_111_192 ();
 FILLCELL_X32 FILLCELL_111_224 ();
 FILLCELL_X32 FILLCELL_111_256 ();
 FILLCELL_X32 FILLCELL_111_288 ();
 FILLCELL_X32 FILLCELL_111_320 ();
 FILLCELL_X32 FILLCELL_111_352 ();
 FILLCELL_X32 FILLCELL_111_384 ();
 FILLCELL_X32 FILLCELL_111_416 ();
 FILLCELL_X32 FILLCELL_111_448 ();
 FILLCELL_X32 FILLCELL_111_480 ();
 FILLCELL_X32 FILLCELL_111_512 ();
 FILLCELL_X8 FILLCELL_111_544 ();
 FILLCELL_X2 FILLCELL_111_552 ();
 FILLCELL_X32 FILLCELL_111_557 ();
 FILLCELL_X32 FILLCELL_111_589 ();
 FILLCELL_X32 FILLCELL_111_621 ();
 FILLCELL_X32 FILLCELL_111_653 ();
 FILLCELL_X32 FILLCELL_111_685 ();
 FILLCELL_X32 FILLCELL_111_717 ();
 FILLCELL_X32 FILLCELL_111_749 ();
 FILLCELL_X32 FILLCELL_111_781 ();
 FILLCELL_X32 FILLCELL_111_813 ();
 FILLCELL_X32 FILLCELL_111_845 ();
 FILLCELL_X32 FILLCELL_111_877 ();
 FILLCELL_X32 FILLCELL_111_909 ();
 FILLCELL_X32 FILLCELL_111_941 ();
 FILLCELL_X32 FILLCELL_111_973 ();
 FILLCELL_X32 FILLCELL_111_1005 ();
 FILLCELL_X32 FILLCELL_111_1037 ();
 FILLCELL_X32 FILLCELL_111_1069 ();
 FILLCELL_X32 FILLCELL_111_1101 ();
 FILLCELL_X32 FILLCELL_111_1133 ();
 FILLCELL_X32 FILLCELL_111_1165 ();
 FILLCELL_X32 FILLCELL_111_1197 ();
 FILLCELL_X32 FILLCELL_111_1229 ();
 FILLCELL_X32 FILLCELL_111_1261 ();
 FILLCELL_X32 FILLCELL_111_1293 ();
 FILLCELL_X32 FILLCELL_111_1325 ();
 FILLCELL_X32 FILLCELL_111_1357 ();
 FILLCELL_X32 FILLCELL_111_1389 ();
 FILLCELL_X32 FILLCELL_111_1421 ();
 FILLCELL_X32 FILLCELL_111_1453 ();
 FILLCELL_X32 FILLCELL_111_1485 ();
 FILLCELL_X32 FILLCELL_111_1517 ();
 FILLCELL_X32 FILLCELL_111_1549 ();
 FILLCELL_X32 FILLCELL_111_1581 ();
 FILLCELL_X32 FILLCELL_111_1613 ();
 FILLCELL_X32 FILLCELL_111_1645 ();
 FILLCELL_X32 FILLCELL_111_1677 ();
 FILLCELL_X32 FILLCELL_111_1709 ();
 FILLCELL_X32 FILLCELL_111_1741 ();
 FILLCELL_X32 FILLCELL_111_1773 ();
 FILLCELL_X32 FILLCELL_111_1805 ();
 FILLCELL_X32 FILLCELL_111_1837 ();
 FILLCELL_X16 FILLCELL_111_1869 ();
 FILLCELL_X8 FILLCELL_111_1885 ();
 FILLCELL_X4 FILLCELL_111_1893 ();
 FILLCELL_X32 FILLCELL_112_0 ();
 FILLCELL_X32 FILLCELL_112_32 ();
 FILLCELL_X32 FILLCELL_112_64 ();
 FILLCELL_X32 FILLCELL_112_96 ();
 FILLCELL_X32 FILLCELL_112_128 ();
 FILLCELL_X32 FILLCELL_112_160 ();
 FILLCELL_X32 FILLCELL_112_192 ();
 FILLCELL_X32 FILLCELL_112_227 ();
 FILLCELL_X32 FILLCELL_112_259 ();
 FILLCELL_X32 FILLCELL_112_291 ();
 FILLCELL_X32 FILLCELL_112_323 ();
 FILLCELL_X32 FILLCELL_112_355 ();
 FILLCELL_X32 FILLCELL_112_387 ();
 FILLCELL_X32 FILLCELL_112_419 ();
 FILLCELL_X32 FILLCELL_112_451 ();
 FILLCELL_X32 FILLCELL_112_483 ();
 FILLCELL_X32 FILLCELL_112_515 ();
 FILLCELL_X16 FILLCELL_112_547 ();
 FILLCELL_X8 FILLCELL_112_563 ();
 FILLCELL_X2 FILLCELL_112_571 ();
 FILLCELL_X32 FILLCELL_112_578 ();
 FILLCELL_X32 FILLCELL_112_610 ();
 FILLCELL_X32 FILLCELL_112_642 ();
 FILLCELL_X32 FILLCELL_112_674 ();
 FILLCELL_X32 FILLCELL_112_706 ();
 FILLCELL_X32 FILLCELL_112_738 ();
 FILLCELL_X32 FILLCELL_112_770 ();
 FILLCELL_X32 FILLCELL_112_802 ();
 FILLCELL_X32 FILLCELL_112_834 ();
 FILLCELL_X32 FILLCELL_112_866 ();
 FILLCELL_X32 FILLCELL_112_898 ();
 FILLCELL_X32 FILLCELL_112_930 ();
 FILLCELL_X32 FILLCELL_112_962 ();
 FILLCELL_X32 FILLCELL_112_994 ();
 FILLCELL_X32 FILLCELL_112_1026 ();
 FILLCELL_X32 FILLCELL_112_1058 ();
 FILLCELL_X32 FILLCELL_112_1090 ();
 FILLCELL_X32 FILLCELL_112_1122 ();
 FILLCELL_X16 FILLCELL_112_1154 ();
 FILLCELL_X8 FILLCELL_112_1170 ();
 FILLCELL_X32 FILLCELL_112_1195 ();
 FILLCELL_X32 FILLCELL_112_1227 ();
 FILLCELL_X32 FILLCELL_112_1259 ();
 FILLCELL_X32 FILLCELL_112_1291 ();
 FILLCELL_X32 FILLCELL_112_1323 ();
 FILLCELL_X32 FILLCELL_112_1355 ();
 FILLCELL_X32 FILLCELL_112_1387 ();
 FILLCELL_X32 FILLCELL_112_1419 ();
 FILLCELL_X32 FILLCELL_112_1451 ();
 FILLCELL_X32 FILLCELL_112_1483 ();
 FILLCELL_X32 FILLCELL_112_1515 ();
 FILLCELL_X32 FILLCELL_112_1547 ();
 FILLCELL_X32 FILLCELL_112_1579 ();
 FILLCELL_X32 FILLCELL_112_1611 ();
 FILLCELL_X32 FILLCELL_112_1643 ();
 FILLCELL_X32 FILLCELL_112_1675 ();
 FILLCELL_X32 FILLCELL_112_1707 ();
 FILLCELL_X32 FILLCELL_112_1739 ();
 FILLCELL_X32 FILLCELL_112_1771 ();
 FILLCELL_X32 FILLCELL_112_1803 ();
 FILLCELL_X32 FILLCELL_112_1835 ();
 FILLCELL_X16 FILLCELL_112_1867 ();
 FILLCELL_X8 FILLCELL_112_1883 ();
 FILLCELL_X4 FILLCELL_112_1891 ();
 FILLCELL_X2 FILLCELL_112_1895 ();
 FILLCELL_X32 FILLCELL_113_0 ();
 FILLCELL_X32 FILLCELL_113_32 ();
 FILLCELL_X32 FILLCELL_113_64 ();
 FILLCELL_X32 FILLCELL_113_96 ();
 FILLCELL_X32 FILLCELL_113_128 ();
 FILLCELL_X32 FILLCELL_113_160 ();
 FILLCELL_X32 FILLCELL_113_192 ();
 FILLCELL_X32 FILLCELL_113_224 ();
 FILLCELL_X32 FILLCELL_113_256 ();
 FILLCELL_X32 FILLCELL_113_288 ();
 FILLCELL_X32 FILLCELL_113_320 ();
 FILLCELL_X32 FILLCELL_113_352 ();
 FILLCELL_X32 FILLCELL_113_384 ();
 FILLCELL_X32 FILLCELL_113_416 ();
 FILLCELL_X32 FILLCELL_113_448 ();
 FILLCELL_X32 FILLCELL_113_480 ();
 FILLCELL_X32 FILLCELL_113_512 ();
 FILLCELL_X16 FILLCELL_113_544 ();
 FILLCELL_X4 FILLCELL_113_560 ();
 FILLCELL_X32 FILLCELL_113_568 ();
 FILLCELL_X32 FILLCELL_113_600 ();
 FILLCELL_X32 FILLCELL_113_632 ();
 FILLCELL_X32 FILLCELL_113_664 ();
 FILLCELL_X32 FILLCELL_113_696 ();
 FILLCELL_X32 FILLCELL_113_728 ();
 FILLCELL_X32 FILLCELL_113_760 ();
 FILLCELL_X32 FILLCELL_113_792 ();
 FILLCELL_X32 FILLCELL_113_824 ();
 FILLCELL_X32 FILLCELL_113_856 ();
 FILLCELL_X32 FILLCELL_113_888 ();
 FILLCELL_X32 FILLCELL_113_920 ();
 FILLCELL_X32 FILLCELL_113_952 ();
 FILLCELL_X32 FILLCELL_113_984 ();
 FILLCELL_X32 FILLCELL_113_1016 ();
 FILLCELL_X32 FILLCELL_113_1048 ();
 FILLCELL_X32 FILLCELL_113_1080 ();
 FILLCELL_X32 FILLCELL_113_1112 ();
 FILLCELL_X16 FILLCELL_113_1144 ();
 FILLCELL_X8 FILLCELL_113_1160 ();
 FILLCELL_X4 FILLCELL_113_1168 ();
 FILLCELL_X2 FILLCELL_113_1172 ();
 FILLCELL_X1 FILLCELL_113_1174 ();
 FILLCELL_X32 FILLCELL_113_1178 ();
 FILLCELL_X32 FILLCELL_113_1210 ();
 FILLCELL_X32 FILLCELL_113_1242 ();
 FILLCELL_X32 FILLCELL_113_1274 ();
 FILLCELL_X32 FILLCELL_113_1306 ();
 FILLCELL_X32 FILLCELL_113_1338 ();
 FILLCELL_X32 FILLCELL_113_1370 ();
 FILLCELL_X32 FILLCELL_113_1402 ();
 FILLCELL_X32 FILLCELL_113_1434 ();
 FILLCELL_X32 FILLCELL_113_1466 ();
 FILLCELL_X32 FILLCELL_113_1498 ();
 FILLCELL_X32 FILLCELL_113_1530 ();
 FILLCELL_X32 FILLCELL_113_1562 ();
 FILLCELL_X32 FILLCELL_113_1594 ();
 FILLCELL_X32 FILLCELL_113_1626 ();
 FILLCELL_X32 FILLCELL_113_1658 ();
 FILLCELL_X32 FILLCELL_113_1690 ();
 FILLCELL_X32 FILLCELL_113_1722 ();
 FILLCELL_X32 FILLCELL_113_1754 ();
 FILLCELL_X32 FILLCELL_113_1786 ();
 FILLCELL_X32 FILLCELL_113_1818 ();
 FILLCELL_X32 FILLCELL_113_1850 ();
 FILLCELL_X8 FILLCELL_113_1882 ();
 FILLCELL_X4 FILLCELL_113_1890 ();
 FILLCELL_X2 FILLCELL_113_1894 ();
 FILLCELL_X1 FILLCELL_113_1896 ();
 FILLCELL_X32 FILLCELL_114_0 ();
 FILLCELL_X32 FILLCELL_114_32 ();
 FILLCELL_X32 FILLCELL_114_64 ();
 FILLCELL_X32 FILLCELL_114_96 ();
 FILLCELL_X32 FILLCELL_114_128 ();
 FILLCELL_X32 FILLCELL_114_160 ();
 FILLCELL_X32 FILLCELL_114_192 ();
 FILLCELL_X32 FILLCELL_114_224 ();
 FILLCELL_X32 FILLCELL_114_256 ();
 FILLCELL_X32 FILLCELL_114_288 ();
 FILLCELL_X32 FILLCELL_114_320 ();
 FILLCELL_X32 FILLCELL_114_352 ();
 FILLCELL_X32 FILLCELL_114_384 ();
 FILLCELL_X32 FILLCELL_114_416 ();
 FILLCELL_X32 FILLCELL_114_448 ();
 FILLCELL_X32 FILLCELL_114_480 ();
 FILLCELL_X32 FILLCELL_114_512 ();
 FILLCELL_X32 FILLCELL_114_544 ();
 FILLCELL_X8 FILLCELL_114_576 ();
 FILLCELL_X2 FILLCELL_114_584 ();
 FILLCELL_X1 FILLCELL_114_586 ();
 FILLCELL_X32 FILLCELL_114_590 ();
 FILLCELL_X32 FILLCELL_114_622 ();
 FILLCELL_X16 FILLCELL_114_654 ();
 FILLCELL_X4 FILLCELL_114_670 ();
 FILLCELL_X2 FILLCELL_114_674 ();
 FILLCELL_X32 FILLCELL_114_679 ();
 FILLCELL_X32 FILLCELL_114_711 ();
 FILLCELL_X32 FILLCELL_114_743 ();
 FILLCELL_X32 FILLCELL_114_775 ();
 FILLCELL_X32 FILLCELL_114_807 ();
 FILLCELL_X16 FILLCELL_114_839 ();
 FILLCELL_X2 FILLCELL_114_855 ();
 FILLCELL_X32 FILLCELL_114_861 ();
 FILLCELL_X16 FILLCELL_114_893 ();
 FILLCELL_X8 FILLCELL_114_909 ();
 FILLCELL_X2 FILLCELL_114_917 ();
 FILLCELL_X32 FILLCELL_114_923 ();
 FILLCELL_X32 FILLCELL_114_955 ();
 FILLCELL_X32 FILLCELL_114_987 ();
 FILLCELL_X32 FILLCELL_114_1019 ();
 FILLCELL_X32 FILLCELL_114_1051 ();
 FILLCELL_X32 FILLCELL_114_1083 ();
 FILLCELL_X32 FILLCELL_114_1115 ();
 FILLCELL_X32 FILLCELL_114_1147 ();
 FILLCELL_X32 FILLCELL_114_1179 ();
 FILLCELL_X32 FILLCELL_114_1211 ();
 FILLCELL_X32 FILLCELL_114_1243 ();
 FILLCELL_X32 FILLCELL_114_1275 ();
 FILLCELL_X32 FILLCELL_114_1307 ();
 FILLCELL_X32 FILLCELL_114_1339 ();
 FILLCELL_X32 FILLCELL_114_1371 ();
 FILLCELL_X32 FILLCELL_114_1403 ();
 FILLCELL_X32 FILLCELL_114_1435 ();
 FILLCELL_X32 FILLCELL_114_1467 ();
 FILLCELL_X32 FILLCELL_114_1499 ();
 FILLCELL_X32 FILLCELL_114_1531 ();
 FILLCELL_X32 FILLCELL_114_1563 ();
 FILLCELL_X32 FILLCELL_114_1595 ();
 FILLCELL_X32 FILLCELL_114_1627 ();
 FILLCELL_X32 FILLCELL_114_1659 ();
 FILLCELL_X32 FILLCELL_114_1691 ();
 FILLCELL_X32 FILLCELL_114_1723 ();
 FILLCELL_X32 FILLCELL_114_1755 ();
 FILLCELL_X32 FILLCELL_114_1787 ();
 FILLCELL_X32 FILLCELL_114_1819 ();
 FILLCELL_X32 FILLCELL_114_1851 ();
 FILLCELL_X8 FILLCELL_114_1883 ();
 FILLCELL_X4 FILLCELL_114_1891 ();
 FILLCELL_X2 FILLCELL_114_1895 ();
 FILLCELL_X32 FILLCELL_115_0 ();
 FILLCELL_X32 FILLCELL_115_32 ();
 FILLCELL_X16 FILLCELL_115_64 ();
 FILLCELL_X4 FILLCELL_115_80 ();
 FILLCELL_X32 FILLCELL_115_87 ();
 FILLCELL_X32 FILLCELL_115_119 ();
 FILLCELL_X32 FILLCELL_115_151 ();
 FILLCELL_X32 FILLCELL_115_183 ();
 FILLCELL_X32 FILLCELL_115_215 ();
 FILLCELL_X32 FILLCELL_115_247 ();
 FILLCELL_X32 FILLCELL_115_279 ();
 FILLCELL_X32 FILLCELL_115_311 ();
 FILLCELL_X32 FILLCELL_115_343 ();
 FILLCELL_X32 FILLCELL_115_375 ();
 FILLCELL_X32 FILLCELL_115_407 ();
 FILLCELL_X2 FILLCELL_115_439 ();
 FILLCELL_X32 FILLCELL_115_445 ();
 FILLCELL_X32 FILLCELL_115_477 ();
 FILLCELL_X32 FILLCELL_115_509 ();
 FILLCELL_X32 FILLCELL_115_541 ();
 FILLCELL_X32 FILLCELL_115_573 ();
 FILLCELL_X32 FILLCELL_115_605 ();
 FILLCELL_X32 FILLCELL_115_637 ();
 FILLCELL_X8 FILLCELL_115_669 ();
 FILLCELL_X2 FILLCELL_115_677 ();
 FILLCELL_X1 FILLCELL_115_679 ();
 FILLCELL_X32 FILLCELL_115_682 ();
 FILLCELL_X32 FILLCELL_115_714 ();
 FILLCELL_X32 FILLCELL_115_746 ();
 FILLCELL_X32 FILLCELL_115_778 ();
 FILLCELL_X32 FILLCELL_115_810 ();
 FILLCELL_X32 FILLCELL_115_842 ();
 FILLCELL_X32 FILLCELL_115_874 ();
 FILLCELL_X32 FILLCELL_115_906 ();
 FILLCELL_X32 FILLCELL_115_938 ();
 FILLCELL_X32 FILLCELL_115_970 ();
 FILLCELL_X32 FILLCELL_115_1002 ();
 FILLCELL_X32 FILLCELL_115_1034 ();
 FILLCELL_X32 FILLCELL_115_1066 ();
 FILLCELL_X32 FILLCELL_115_1098 ();
 FILLCELL_X32 FILLCELL_115_1130 ();
 FILLCELL_X32 FILLCELL_115_1162 ();
 FILLCELL_X32 FILLCELL_115_1194 ();
 FILLCELL_X32 FILLCELL_115_1226 ();
 FILLCELL_X32 FILLCELL_115_1258 ();
 FILLCELL_X32 FILLCELL_115_1290 ();
 FILLCELL_X32 FILLCELL_115_1322 ();
 FILLCELL_X32 FILLCELL_115_1354 ();
 FILLCELL_X32 FILLCELL_115_1386 ();
 FILLCELL_X32 FILLCELL_115_1418 ();
 FILLCELL_X32 FILLCELL_115_1450 ();
 FILLCELL_X32 FILLCELL_115_1482 ();
 FILLCELL_X32 FILLCELL_115_1514 ();
 FILLCELL_X32 FILLCELL_115_1546 ();
 FILLCELL_X32 FILLCELL_115_1578 ();
 FILLCELL_X32 FILLCELL_115_1610 ();
 FILLCELL_X32 FILLCELL_115_1642 ();
 FILLCELL_X32 FILLCELL_115_1674 ();
 FILLCELL_X32 FILLCELL_115_1706 ();
 FILLCELL_X32 FILLCELL_115_1738 ();
 FILLCELL_X32 FILLCELL_115_1770 ();
 FILLCELL_X32 FILLCELL_115_1802 ();
 FILLCELL_X32 FILLCELL_115_1834 ();
 FILLCELL_X16 FILLCELL_115_1866 ();
 FILLCELL_X8 FILLCELL_115_1882 ();
 FILLCELL_X4 FILLCELL_115_1890 ();
 FILLCELL_X2 FILLCELL_115_1894 ();
 FILLCELL_X1 FILLCELL_115_1896 ();
 FILLCELL_X32 FILLCELL_116_0 ();
 FILLCELL_X32 FILLCELL_116_32 ();
 FILLCELL_X32 FILLCELL_116_64 ();
 FILLCELL_X32 FILLCELL_116_96 ();
 FILLCELL_X32 FILLCELL_116_128 ();
 FILLCELL_X32 FILLCELL_116_160 ();
 FILLCELL_X32 FILLCELL_116_192 ();
 FILLCELL_X32 FILLCELL_116_224 ();
 FILLCELL_X32 FILLCELL_116_256 ();
 FILLCELL_X32 FILLCELL_116_288 ();
 FILLCELL_X32 FILLCELL_116_320 ();
 FILLCELL_X32 FILLCELL_116_352 ();
 FILLCELL_X32 FILLCELL_116_384 ();
 FILLCELL_X32 FILLCELL_116_416 ();
 FILLCELL_X32 FILLCELL_116_448 ();
 FILLCELL_X32 FILLCELL_116_480 ();
 FILLCELL_X32 FILLCELL_116_512 ();
 FILLCELL_X8 FILLCELL_116_544 ();
 FILLCELL_X1 FILLCELL_116_552 ();
 FILLCELL_X32 FILLCELL_116_555 ();
 FILLCELL_X32 FILLCELL_116_587 ();
 FILLCELL_X32 FILLCELL_116_619 ();
 FILLCELL_X32 FILLCELL_116_651 ();
 FILLCELL_X32 FILLCELL_116_683 ();
 FILLCELL_X32 FILLCELL_116_715 ();
 FILLCELL_X32 FILLCELL_116_747 ();
 FILLCELL_X32 FILLCELL_116_779 ();
 FILLCELL_X16 FILLCELL_116_811 ();
 FILLCELL_X4 FILLCELL_116_827 ();
 FILLCELL_X2 FILLCELL_116_831 ();
 FILLCELL_X1 FILLCELL_116_833 ();
 FILLCELL_X32 FILLCELL_116_839 ();
 FILLCELL_X32 FILLCELL_116_871 ();
 FILLCELL_X32 FILLCELL_116_903 ();
 FILLCELL_X16 FILLCELL_116_935 ();
 FILLCELL_X4 FILLCELL_116_951 ();
 FILLCELL_X2 FILLCELL_116_955 ();
 FILLCELL_X32 FILLCELL_116_960 ();
 FILLCELL_X32 FILLCELL_116_992 ();
 FILLCELL_X32 FILLCELL_116_1024 ();
 FILLCELL_X32 FILLCELL_116_1056 ();
 FILLCELL_X32 FILLCELL_116_1088 ();
 FILLCELL_X32 FILLCELL_116_1120 ();
 FILLCELL_X32 FILLCELL_116_1152 ();
 FILLCELL_X32 FILLCELL_116_1184 ();
 FILLCELL_X32 FILLCELL_116_1216 ();
 FILLCELL_X32 FILLCELL_116_1248 ();
 FILLCELL_X32 FILLCELL_116_1280 ();
 FILLCELL_X32 FILLCELL_116_1312 ();
 FILLCELL_X32 FILLCELL_116_1344 ();
 FILLCELL_X32 FILLCELL_116_1376 ();
 FILLCELL_X32 FILLCELL_116_1408 ();
 FILLCELL_X32 FILLCELL_116_1440 ();
 FILLCELL_X32 FILLCELL_116_1472 ();
 FILLCELL_X32 FILLCELL_116_1504 ();
 FILLCELL_X32 FILLCELL_116_1536 ();
 FILLCELL_X32 FILLCELL_116_1568 ();
 FILLCELL_X32 FILLCELL_116_1600 ();
 FILLCELL_X32 FILLCELL_116_1632 ();
 FILLCELL_X32 FILLCELL_116_1664 ();
 FILLCELL_X32 FILLCELL_116_1696 ();
 FILLCELL_X32 FILLCELL_116_1728 ();
 FILLCELL_X32 FILLCELL_116_1760 ();
 FILLCELL_X32 FILLCELL_116_1792 ();
 FILLCELL_X32 FILLCELL_116_1824 ();
 FILLCELL_X32 FILLCELL_116_1856 ();
 FILLCELL_X8 FILLCELL_116_1888 ();
 FILLCELL_X1 FILLCELL_116_1896 ();
 FILLCELL_X32 FILLCELL_117_0 ();
 FILLCELL_X4 FILLCELL_117_32 ();
 FILLCELL_X1 FILLCELL_117_36 ();
 FILLCELL_X32 FILLCELL_117_54 ();
 FILLCELL_X16 FILLCELL_117_86 ();
 FILLCELL_X4 FILLCELL_117_102 ();
 FILLCELL_X32 FILLCELL_117_110 ();
 FILLCELL_X32 FILLCELL_117_142 ();
 FILLCELL_X32 FILLCELL_117_174 ();
 FILLCELL_X32 FILLCELL_117_206 ();
 FILLCELL_X32 FILLCELL_117_238 ();
 FILLCELL_X32 FILLCELL_117_270 ();
 FILLCELL_X32 FILLCELL_117_302 ();
 FILLCELL_X32 FILLCELL_117_334 ();
 FILLCELL_X32 FILLCELL_117_366 ();
 FILLCELL_X32 FILLCELL_117_398 ();
 FILLCELL_X32 FILLCELL_117_430 ();
 FILLCELL_X8 FILLCELL_117_462 ();
 FILLCELL_X32 FILLCELL_117_479 ();
 FILLCELL_X32 FILLCELL_117_511 ();
 FILLCELL_X32 FILLCELL_117_543 ();
 FILLCELL_X32 FILLCELL_117_575 ();
 FILLCELL_X32 FILLCELL_117_607 ();
 FILLCELL_X32 FILLCELL_117_639 ();
 FILLCELL_X32 FILLCELL_117_671 ();
 FILLCELL_X32 FILLCELL_117_703 ();
 FILLCELL_X32 FILLCELL_117_735 ();
 FILLCELL_X32 FILLCELL_117_767 ();
 FILLCELL_X32 FILLCELL_117_799 ();
 FILLCELL_X32 FILLCELL_117_831 ();
 FILLCELL_X8 FILLCELL_117_863 ();
 FILLCELL_X1 FILLCELL_117_871 ();
 FILLCELL_X32 FILLCELL_117_876 ();
 FILLCELL_X8 FILLCELL_117_908 ();
 FILLCELL_X2 FILLCELL_117_916 ();
 FILLCELL_X8 FILLCELL_117_922 ();
 FILLCELL_X2 FILLCELL_117_930 ();
 FILLCELL_X1 FILLCELL_117_932 ();
 FILLCELL_X32 FILLCELL_117_937 ();
 FILLCELL_X16 FILLCELL_117_969 ();
 FILLCELL_X8 FILLCELL_117_985 ();
 FILLCELL_X4 FILLCELL_117_993 ();
 FILLCELL_X1 FILLCELL_117_997 ();
 FILLCELL_X32 FILLCELL_117_1001 ();
 FILLCELL_X32 FILLCELL_117_1033 ();
 FILLCELL_X8 FILLCELL_117_1065 ();
 FILLCELL_X32 FILLCELL_117_1090 ();
 FILLCELL_X32 FILLCELL_117_1122 ();
 FILLCELL_X32 FILLCELL_117_1154 ();
 FILLCELL_X32 FILLCELL_117_1186 ();
 FILLCELL_X32 FILLCELL_117_1218 ();
 FILLCELL_X32 FILLCELL_117_1250 ();
 FILLCELL_X32 FILLCELL_117_1282 ();
 FILLCELL_X32 FILLCELL_117_1314 ();
 FILLCELL_X32 FILLCELL_117_1346 ();
 FILLCELL_X32 FILLCELL_117_1378 ();
 FILLCELL_X32 FILLCELL_117_1410 ();
 FILLCELL_X32 FILLCELL_117_1442 ();
 FILLCELL_X32 FILLCELL_117_1474 ();
 FILLCELL_X32 FILLCELL_117_1506 ();
 FILLCELL_X32 FILLCELL_117_1538 ();
 FILLCELL_X32 FILLCELL_117_1570 ();
 FILLCELL_X32 FILLCELL_117_1602 ();
 FILLCELL_X32 FILLCELL_117_1634 ();
 FILLCELL_X32 FILLCELL_117_1666 ();
 FILLCELL_X32 FILLCELL_117_1698 ();
 FILLCELL_X32 FILLCELL_117_1730 ();
 FILLCELL_X32 FILLCELL_117_1762 ();
 FILLCELL_X32 FILLCELL_117_1794 ();
 FILLCELL_X32 FILLCELL_117_1826 ();
 FILLCELL_X32 FILLCELL_117_1858 ();
 FILLCELL_X4 FILLCELL_117_1890 ();
 FILLCELL_X2 FILLCELL_117_1894 ();
 FILLCELL_X1 FILLCELL_117_1896 ();
 FILLCELL_X32 FILLCELL_118_0 ();
 FILLCELL_X32 FILLCELL_118_32 ();
 FILLCELL_X16 FILLCELL_118_64 ();
 FILLCELL_X8 FILLCELL_118_80 ();
 FILLCELL_X32 FILLCELL_118_92 ();
 FILLCELL_X32 FILLCELL_118_124 ();
 FILLCELL_X16 FILLCELL_118_156 ();
 FILLCELL_X8 FILLCELL_118_172 ();
 FILLCELL_X4 FILLCELL_118_180 ();
 FILLCELL_X4 FILLCELL_118_201 ();
 FILLCELL_X32 FILLCELL_118_209 ();
 FILLCELL_X32 FILLCELL_118_241 ();
 FILLCELL_X32 FILLCELL_118_273 ();
 FILLCELL_X32 FILLCELL_118_305 ();
 FILLCELL_X32 FILLCELL_118_337 ();
 FILLCELL_X8 FILLCELL_118_369 ();
 FILLCELL_X1 FILLCELL_118_377 ();
 FILLCELL_X4 FILLCELL_118_381 ();
 FILLCELL_X2 FILLCELL_118_385 ();
 FILLCELL_X1 FILLCELL_118_387 ();
 FILLCELL_X32 FILLCELL_118_390 ();
 FILLCELL_X16 FILLCELL_118_422 ();
 FILLCELL_X4 FILLCELL_118_438 ();
 FILLCELL_X32 FILLCELL_118_444 ();
 FILLCELL_X32 FILLCELL_118_476 ();
 FILLCELL_X16 FILLCELL_118_508 ();
 FILLCELL_X8 FILLCELL_118_524 ();
 FILLCELL_X2 FILLCELL_118_532 ();
 FILLCELL_X32 FILLCELL_118_538 ();
 FILLCELL_X32 FILLCELL_118_570 ();
 FILLCELL_X32 FILLCELL_118_602 ();
 FILLCELL_X16 FILLCELL_118_634 ();
 FILLCELL_X8 FILLCELL_118_650 ();
 FILLCELL_X4 FILLCELL_118_658 ();
 FILLCELL_X1 FILLCELL_118_662 ();
 FILLCELL_X8 FILLCELL_118_665 ();
 FILLCELL_X4 FILLCELL_118_673 ();
 FILLCELL_X32 FILLCELL_118_682 ();
 FILLCELL_X32 FILLCELL_118_714 ();
 FILLCELL_X32 FILLCELL_118_746 ();
 FILLCELL_X32 FILLCELL_118_778 ();
 FILLCELL_X32 FILLCELL_118_810 ();
 FILLCELL_X32 FILLCELL_118_842 ();
 FILLCELL_X32 FILLCELL_118_874 ();
 FILLCELL_X32 FILLCELL_118_906 ();
 FILLCELL_X32 FILLCELL_118_938 ();
 FILLCELL_X32 FILLCELL_118_970 ();
 FILLCELL_X8 FILLCELL_118_1002 ();
 FILLCELL_X2 FILLCELL_118_1010 ();
 FILLCELL_X1 FILLCELL_118_1012 ();
 FILLCELL_X32 FILLCELL_118_1017 ();
 FILLCELL_X32 FILLCELL_118_1049 ();
 FILLCELL_X32 FILLCELL_118_1081 ();
 FILLCELL_X32 FILLCELL_118_1113 ();
 FILLCELL_X32 FILLCELL_118_1145 ();
 FILLCELL_X32 FILLCELL_118_1177 ();
 FILLCELL_X32 FILLCELL_118_1209 ();
 FILLCELL_X32 FILLCELL_118_1241 ();
 FILLCELL_X32 FILLCELL_118_1273 ();
 FILLCELL_X32 FILLCELL_118_1305 ();
 FILLCELL_X32 FILLCELL_118_1337 ();
 FILLCELL_X32 FILLCELL_118_1369 ();
 FILLCELL_X32 FILLCELL_118_1401 ();
 FILLCELL_X32 FILLCELL_118_1433 ();
 FILLCELL_X32 FILLCELL_118_1465 ();
 FILLCELL_X32 FILLCELL_118_1497 ();
 FILLCELL_X32 FILLCELL_118_1529 ();
 FILLCELL_X32 FILLCELL_118_1561 ();
 FILLCELL_X32 FILLCELL_118_1593 ();
 FILLCELL_X32 FILLCELL_118_1625 ();
 FILLCELL_X32 FILLCELL_118_1657 ();
 FILLCELL_X32 FILLCELL_118_1689 ();
 FILLCELL_X32 FILLCELL_118_1721 ();
 FILLCELL_X32 FILLCELL_118_1753 ();
 FILLCELL_X32 FILLCELL_118_1785 ();
 FILLCELL_X32 FILLCELL_118_1817 ();
 FILLCELL_X32 FILLCELL_118_1849 ();
 FILLCELL_X16 FILLCELL_118_1881 ();
 FILLCELL_X32 FILLCELL_119_0 ();
 FILLCELL_X32 FILLCELL_119_32 ();
 FILLCELL_X32 FILLCELL_119_64 ();
 FILLCELL_X32 FILLCELL_119_96 ();
 FILLCELL_X32 FILLCELL_119_128 ();
 FILLCELL_X32 FILLCELL_119_160 ();
 FILLCELL_X32 FILLCELL_119_192 ();
 FILLCELL_X32 FILLCELL_119_224 ();
 FILLCELL_X32 FILLCELL_119_256 ();
 FILLCELL_X32 FILLCELL_119_288 ();
 FILLCELL_X8 FILLCELL_119_320 ();
 FILLCELL_X2 FILLCELL_119_328 ();
 FILLCELL_X32 FILLCELL_119_333 ();
 FILLCELL_X32 FILLCELL_119_365 ();
 FILLCELL_X32 FILLCELL_119_397 ();
 FILLCELL_X32 FILLCELL_119_429 ();
 FILLCELL_X32 FILLCELL_119_461 ();
 FILLCELL_X32 FILLCELL_119_493 ();
 FILLCELL_X32 FILLCELL_119_525 ();
 FILLCELL_X16 FILLCELL_119_557 ();
 FILLCELL_X1 FILLCELL_119_573 ();
 FILLCELL_X32 FILLCELL_119_577 ();
 FILLCELL_X32 FILLCELL_119_609 ();
 FILLCELL_X8 FILLCELL_119_641 ();
 FILLCELL_X4 FILLCELL_119_649 ();
 FILLCELL_X2 FILLCELL_119_653 ();
 FILLCELL_X32 FILLCELL_119_660 ();
 FILLCELL_X32 FILLCELL_119_692 ();
 FILLCELL_X32 FILLCELL_119_724 ();
 FILLCELL_X32 FILLCELL_119_756 ();
 FILLCELL_X4 FILLCELL_119_788 ();
 FILLCELL_X2 FILLCELL_119_792 ();
 FILLCELL_X32 FILLCELL_119_797 ();
 FILLCELL_X32 FILLCELL_119_829 ();
 FILLCELL_X32 FILLCELL_119_861 ();
 FILLCELL_X32 FILLCELL_119_893 ();
 FILLCELL_X32 FILLCELL_119_925 ();
 FILLCELL_X32 FILLCELL_119_957 ();
 FILLCELL_X8 FILLCELL_119_989 ();
 FILLCELL_X4 FILLCELL_119_997 ();
 FILLCELL_X2 FILLCELL_119_1001 ();
 FILLCELL_X2 FILLCELL_119_1007 ();
 FILLCELL_X1 FILLCELL_119_1009 ();
 FILLCELL_X32 FILLCELL_119_1013 ();
 FILLCELL_X32 FILLCELL_119_1045 ();
 FILLCELL_X32 FILLCELL_119_1077 ();
 FILLCELL_X32 FILLCELL_119_1109 ();
 FILLCELL_X32 FILLCELL_119_1141 ();
 FILLCELL_X32 FILLCELL_119_1173 ();
 FILLCELL_X32 FILLCELL_119_1205 ();
 FILLCELL_X32 FILLCELL_119_1237 ();
 FILLCELL_X32 FILLCELL_119_1269 ();
 FILLCELL_X32 FILLCELL_119_1301 ();
 FILLCELL_X32 FILLCELL_119_1333 ();
 FILLCELL_X32 FILLCELL_119_1365 ();
 FILLCELL_X32 FILLCELL_119_1397 ();
 FILLCELL_X32 FILLCELL_119_1429 ();
 FILLCELL_X32 FILLCELL_119_1461 ();
 FILLCELL_X32 FILLCELL_119_1493 ();
 FILLCELL_X32 FILLCELL_119_1525 ();
 FILLCELL_X32 FILLCELL_119_1557 ();
 FILLCELL_X32 FILLCELL_119_1589 ();
 FILLCELL_X32 FILLCELL_119_1621 ();
 FILLCELL_X32 FILLCELL_119_1653 ();
 FILLCELL_X32 FILLCELL_119_1685 ();
 FILLCELL_X32 FILLCELL_119_1717 ();
 FILLCELL_X32 FILLCELL_119_1749 ();
 FILLCELL_X32 FILLCELL_119_1781 ();
 FILLCELL_X32 FILLCELL_119_1813 ();
 FILLCELL_X32 FILLCELL_119_1845 ();
 FILLCELL_X16 FILLCELL_119_1877 ();
 FILLCELL_X4 FILLCELL_119_1893 ();
 FILLCELL_X32 FILLCELL_120_0 ();
 FILLCELL_X32 FILLCELL_120_32 ();
 FILLCELL_X32 FILLCELL_120_64 ();
 FILLCELL_X32 FILLCELL_120_96 ();
 FILLCELL_X32 FILLCELL_120_128 ();
 FILLCELL_X32 FILLCELL_120_160 ();
 FILLCELL_X32 FILLCELL_120_192 ();
 FILLCELL_X32 FILLCELL_120_224 ();
 FILLCELL_X32 FILLCELL_120_256 ();
 FILLCELL_X32 FILLCELL_120_288 ();
 FILLCELL_X32 FILLCELL_120_320 ();
 FILLCELL_X16 FILLCELL_120_352 ();
 FILLCELL_X32 FILLCELL_120_371 ();
 FILLCELL_X32 FILLCELL_120_403 ();
 FILLCELL_X32 FILLCELL_120_441 ();
 FILLCELL_X32 FILLCELL_120_473 ();
 FILLCELL_X32 FILLCELL_120_505 ();
 FILLCELL_X16 FILLCELL_120_537 ();
 FILLCELL_X8 FILLCELL_120_553 ();
 FILLCELL_X4 FILLCELL_120_561 ();
 FILLCELL_X1 FILLCELL_120_565 ();
 FILLCELL_X32 FILLCELL_120_568 ();
 FILLCELL_X32 FILLCELL_120_600 ();
 FILLCELL_X32 FILLCELL_120_632 ();
 FILLCELL_X32 FILLCELL_120_664 ();
 FILLCELL_X32 FILLCELL_120_696 ();
 FILLCELL_X16 FILLCELL_120_728 ();
 FILLCELL_X1 FILLCELL_120_744 ();
 FILLCELL_X32 FILLCELL_120_750 ();
 FILLCELL_X8 FILLCELL_120_782 ();
 FILLCELL_X2 FILLCELL_120_790 ();
 FILLCELL_X1 FILLCELL_120_792 ();
 FILLCELL_X16 FILLCELL_120_796 ();
 FILLCELL_X32 FILLCELL_120_816 ();
 FILLCELL_X8 FILLCELL_120_848 ();
 FILLCELL_X4 FILLCELL_120_856 ();
 FILLCELL_X1 FILLCELL_120_860 ();
 FILLCELL_X32 FILLCELL_120_867 ();
 FILLCELL_X32 FILLCELL_120_899 ();
 FILLCELL_X32 FILLCELL_120_931 ();
 FILLCELL_X32 FILLCELL_120_963 ();
 FILLCELL_X32 FILLCELL_120_995 ();
 FILLCELL_X32 FILLCELL_120_1027 ();
 FILLCELL_X32 FILLCELL_120_1059 ();
 FILLCELL_X32 FILLCELL_120_1091 ();
 FILLCELL_X32 FILLCELL_120_1123 ();
 FILLCELL_X32 FILLCELL_120_1155 ();
 FILLCELL_X32 FILLCELL_120_1187 ();
 FILLCELL_X32 FILLCELL_120_1219 ();
 FILLCELL_X32 FILLCELL_120_1251 ();
 FILLCELL_X32 FILLCELL_120_1283 ();
 FILLCELL_X32 FILLCELL_120_1315 ();
 FILLCELL_X32 FILLCELL_120_1347 ();
 FILLCELL_X32 FILLCELL_120_1379 ();
 FILLCELL_X32 FILLCELL_120_1411 ();
 FILLCELL_X32 FILLCELL_120_1443 ();
 FILLCELL_X32 FILLCELL_120_1475 ();
 FILLCELL_X32 FILLCELL_120_1507 ();
 FILLCELL_X32 FILLCELL_120_1539 ();
 FILLCELL_X32 FILLCELL_120_1571 ();
 FILLCELL_X32 FILLCELL_120_1603 ();
 FILLCELL_X32 FILLCELL_120_1635 ();
 FILLCELL_X32 FILLCELL_120_1667 ();
 FILLCELL_X32 FILLCELL_120_1699 ();
 FILLCELL_X32 FILLCELL_120_1731 ();
 FILLCELL_X32 FILLCELL_120_1763 ();
 FILLCELL_X32 FILLCELL_120_1795 ();
 FILLCELL_X32 FILLCELL_120_1827 ();
 FILLCELL_X32 FILLCELL_120_1859 ();
 FILLCELL_X4 FILLCELL_120_1891 ();
 FILLCELL_X2 FILLCELL_120_1895 ();
 FILLCELL_X32 FILLCELL_121_0 ();
 FILLCELL_X32 FILLCELL_121_32 ();
 FILLCELL_X32 FILLCELL_121_64 ();
 FILLCELL_X32 FILLCELL_121_96 ();
 FILLCELL_X32 FILLCELL_121_128 ();
 FILLCELL_X32 FILLCELL_121_160 ();
 FILLCELL_X32 FILLCELL_121_192 ();
 FILLCELL_X32 FILLCELL_121_224 ();
 FILLCELL_X32 FILLCELL_121_256 ();
 FILLCELL_X16 FILLCELL_121_288 ();
 FILLCELL_X8 FILLCELL_121_304 ();
 FILLCELL_X4 FILLCELL_121_312 ();
 FILLCELL_X2 FILLCELL_121_316 ();
 FILLCELL_X32 FILLCELL_121_324 ();
 FILLCELL_X32 FILLCELL_121_356 ();
 FILLCELL_X32 FILLCELL_121_388 ();
 FILLCELL_X32 FILLCELL_121_420 ();
 FILLCELL_X32 FILLCELL_121_452 ();
 FILLCELL_X32 FILLCELL_121_484 ();
 FILLCELL_X32 FILLCELL_121_516 ();
 FILLCELL_X32 FILLCELL_121_548 ();
 FILLCELL_X32 FILLCELL_121_580 ();
 FILLCELL_X32 FILLCELL_121_612 ();
 FILLCELL_X8 FILLCELL_121_644 ();
 FILLCELL_X32 FILLCELL_121_656 ();
 FILLCELL_X32 FILLCELL_121_688 ();
 FILLCELL_X16 FILLCELL_121_720 ();
 FILLCELL_X2 FILLCELL_121_736 ();
 FILLCELL_X1 FILLCELL_121_738 ();
 FILLCELL_X32 FILLCELL_121_744 ();
 FILLCELL_X32 FILLCELL_121_776 ();
 FILLCELL_X32 FILLCELL_121_808 ();
 FILLCELL_X32 FILLCELL_121_840 ();
 FILLCELL_X32 FILLCELL_121_872 ();
 FILLCELL_X32 FILLCELL_121_904 ();
 FILLCELL_X32 FILLCELL_121_936 ();
 FILLCELL_X32 FILLCELL_121_968 ();
 FILLCELL_X32 FILLCELL_121_1000 ();
 FILLCELL_X32 FILLCELL_121_1032 ();
 FILLCELL_X32 FILLCELL_121_1064 ();
 FILLCELL_X32 FILLCELL_121_1096 ();
 FILLCELL_X32 FILLCELL_121_1128 ();
 FILLCELL_X32 FILLCELL_121_1160 ();
 FILLCELL_X32 FILLCELL_121_1192 ();
 FILLCELL_X32 FILLCELL_121_1224 ();
 FILLCELL_X32 FILLCELL_121_1256 ();
 FILLCELL_X32 FILLCELL_121_1288 ();
 FILLCELL_X32 FILLCELL_121_1320 ();
 FILLCELL_X32 FILLCELL_121_1352 ();
 FILLCELL_X32 FILLCELL_121_1384 ();
 FILLCELL_X32 FILLCELL_121_1416 ();
 FILLCELL_X32 FILLCELL_121_1448 ();
 FILLCELL_X32 FILLCELL_121_1480 ();
 FILLCELL_X32 FILLCELL_121_1512 ();
 FILLCELL_X32 FILLCELL_121_1544 ();
 FILLCELL_X32 FILLCELL_121_1576 ();
 FILLCELL_X32 FILLCELL_121_1608 ();
 FILLCELL_X32 FILLCELL_121_1640 ();
 FILLCELL_X32 FILLCELL_121_1672 ();
 FILLCELL_X32 FILLCELL_121_1704 ();
 FILLCELL_X32 FILLCELL_121_1736 ();
 FILLCELL_X32 FILLCELL_121_1768 ();
 FILLCELL_X32 FILLCELL_121_1800 ();
 FILLCELL_X32 FILLCELL_121_1832 ();
 FILLCELL_X32 FILLCELL_121_1864 ();
 FILLCELL_X1 FILLCELL_121_1896 ();
 FILLCELL_X32 FILLCELL_122_0 ();
 FILLCELL_X32 FILLCELL_122_32 ();
 FILLCELL_X32 FILLCELL_122_64 ();
 FILLCELL_X32 FILLCELL_122_96 ();
 FILLCELL_X32 FILLCELL_122_128 ();
 FILLCELL_X32 FILLCELL_122_160 ();
 FILLCELL_X32 FILLCELL_122_192 ();
 FILLCELL_X32 FILLCELL_122_224 ();
 FILLCELL_X32 FILLCELL_122_256 ();
 FILLCELL_X32 FILLCELL_122_288 ();
 FILLCELL_X32 FILLCELL_122_320 ();
 FILLCELL_X32 FILLCELL_122_352 ();
 FILLCELL_X32 FILLCELL_122_384 ();
 FILLCELL_X32 FILLCELL_122_416 ();
 FILLCELL_X32 FILLCELL_122_448 ();
 FILLCELL_X32 FILLCELL_122_480 ();
 FILLCELL_X32 FILLCELL_122_512 ();
 FILLCELL_X32 FILLCELL_122_544 ();
 FILLCELL_X32 FILLCELL_122_576 ();
 FILLCELL_X32 FILLCELL_122_608 ();
 FILLCELL_X32 FILLCELL_122_640 ();
 FILLCELL_X32 FILLCELL_122_672 ();
 FILLCELL_X32 FILLCELL_122_704 ();
 FILLCELL_X32 FILLCELL_122_736 ();
 FILLCELL_X32 FILLCELL_122_768 ();
 FILLCELL_X32 FILLCELL_122_800 ();
 FILLCELL_X32 FILLCELL_122_832 ();
 FILLCELL_X32 FILLCELL_122_864 ();
 FILLCELL_X32 FILLCELL_122_896 ();
 FILLCELL_X32 FILLCELL_122_928 ();
 FILLCELL_X32 FILLCELL_122_960 ();
 FILLCELL_X32 FILLCELL_122_992 ();
 FILLCELL_X32 FILLCELL_122_1024 ();
 FILLCELL_X32 FILLCELL_122_1056 ();
 FILLCELL_X32 FILLCELL_122_1088 ();
 FILLCELL_X32 FILLCELL_122_1120 ();
 FILLCELL_X32 FILLCELL_122_1152 ();
 FILLCELL_X32 FILLCELL_122_1184 ();
 FILLCELL_X32 FILLCELL_122_1216 ();
 FILLCELL_X32 FILLCELL_122_1248 ();
 FILLCELL_X32 FILLCELL_122_1280 ();
 FILLCELL_X32 FILLCELL_122_1312 ();
 FILLCELL_X32 FILLCELL_122_1344 ();
 FILLCELL_X32 FILLCELL_122_1376 ();
 FILLCELL_X32 FILLCELL_122_1408 ();
 FILLCELL_X32 FILLCELL_122_1440 ();
 FILLCELL_X32 FILLCELL_122_1472 ();
 FILLCELL_X32 FILLCELL_122_1504 ();
 FILLCELL_X32 FILLCELL_122_1536 ();
 FILLCELL_X32 FILLCELL_122_1568 ();
 FILLCELL_X32 FILLCELL_122_1600 ();
 FILLCELL_X32 FILLCELL_122_1632 ();
 FILLCELL_X32 FILLCELL_122_1664 ();
 FILLCELL_X32 FILLCELL_122_1696 ();
 FILLCELL_X32 FILLCELL_122_1728 ();
 FILLCELL_X32 FILLCELL_122_1760 ();
 FILLCELL_X32 FILLCELL_122_1792 ();
 FILLCELL_X32 FILLCELL_122_1824 ();
 FILLCELL_X32 FILLCELL_122_1856 ();
 FILLCELL_X8 FILLCELL_122_1888 ();
 FILLCELL_X1 FILLCELL_122_1896 ();
 FILLCELL_X32 FILLCELL_123_0 ();
 FILLCELL_X32 FILLCELL_123_32 ();
 FILLCELL_X32 FILLCELL_123_64 ();
 FILLCELL_X32 FILLCELL_123_96 ();
 FILLCELL_X32 FILLCELL_123_128 ();
 FILLCELL_X32 FILLCELL_123_160 ();
 FILLCELL_X32 FILLCELL_123_192 ();
 FILLCELL_X32 FILLCELL_123_224 ();
 FILLCELL_X32 FILLCELL_123_256 ();
 FILLCELL_X8 FILLCELL_123_288 ();
 FILLCELL_X2 FILLCELL_123_296 ();
 FILLCELL_X1 FILLCELL_123_298 ();
 FILLCELL_X32 FILLCELL_123_304 ();
 FILLCELL_X32 FILLCELL_123_336 ();
 FILLCELL_X32 FILLCELL_123_368 ();
 FILLCELL_X32 FILLCELL_123_400 ();
 FILLCELL_X32 FILLCELL_123_432 ();
 FILLCELL_X32 FILLCELL_123_464 ();
 FILLCELL_X32 FILLCELL_123_496 ();
 FILLCELL_X32 FILLCELL_123_528 ();
 FILLCELL_X32 FILLCELL_123_560 ();
 FILLCELL_X32 FILLCELL_123_592 ();
 FILLCELL_X32 FILLCELL_123_624 ();
 FILLCELL_X32 FILLCELL_123_656 ();
 FILLCELL_X32 FILLCELL_123_688 ();
 FILLCELL_X32 FILLCELL_123_720 ();
 FILLCELL_X32 FILLCELL_123_752 ();
 FILLCELL_X32 FILLCELL_123_784 ();
 FILLCELL_X32 FILLCELL_123_816 ();
 FILLCELL_X32 FILLCELL_123_848 ();
 FILLCELL_X32 FILLCELL_123_880 ();
 FILLCELL_X32 FILLCELL_123_912 ();
 FILLCELL_X32 FILLCELL_123_944 ();
 FILLCELL_X32 FILLCELL_123_976 ();
 FILLCELL_X32 FILLCELL_123_1008 ();
 FILLCELL_X32 FILLCELL_123_1040 ();
 FILLCELL_X32 FILLCELL_123_1072 ();
 FILLCELL_X32 FILLCELL_123_1104 ();
 FILLCELL_X32 FILLCELL_123_1136 ();
 FILLCELL_X32 FILLCELL_123_1168 ();
 FILLCELL_X32 FILLCELL_123_1200 ();
 FILLCELL_X32 FILLCELL_123_1232 ();
 FILLCELL_X32 FILLCELL_123_1264 ();
 FILLCELL_X32 FILLCELL_123_1296 ();
 FILLCELL_X32 FILLCELL_123_1328 ();
 FILLCELL_X32 FILLCELL_123_1360 ();
 FILLCELL_X32 FILLCELL_123_1392 ();
 FILLCELL_X32 FILLCELL_123_1424 ();
 FILLCELL_X32 FILLCELL_123_1456 ();
 FILLCELL_X32 FILLCELL_123_1488 ();
 FILLCELL_X32 FILLCELL_123_1520 ();
 FILLCELL_X32 FILLCELL_123_1552 ();
 FILLCELL_X32 FILLCELL_123_1584 ();
 FILLCELL_X32 FILLCELL_123_1616 ();
 FILLCELL_X32 FILLCELL_123_1648 ();
 FILLCELL_X32 FILLCELL_123_1680 ();
 FILLCELL_X32 FILLCELL_123_1712 ();
 FILLCELL_X32 FILLCELL_123_1744 ();
 FILLCELL_X32 FILLCELL_123_1776 ();
 FILLCELL_X32 FILLCELL_123_1808 ();
 FILLCELL_X32 FILLCELL_123_1840 ();
 FILLCELL_X16 FILLCELL_123_1872 ();
 FILLCELL_X8 FILLCELL_123_1888 ();
 FILLCELL_X1 FILLCELL_123_1896 ();
 FILLCELL_X32 FILLCELL_124_0 ();
 FILLCELL_X32 FILLCELL_124_32 ();
 FILLCELL_X32 FILLCELL_124_64 ();
 FILLCELL_X32 FILLCELL_124_96 ();
 FILLCELL_X32 FILLCELL_124_128 ();
 FILLCELL_X16 FILLCELL_124_160 ();
 FILLCELL_X8 FILLCELL_124_176 ();
 FILLCELL_X4 FILLCELL_124_184 ();
 FILLCELL_X1 FILLCELL_124_188 ();
 FILLCELL_X32 FILLCELL_124_192 ();
 FILLCELL_X32 FILLCELL_124_224 ();
 FILLCELL_X32 FILLCELL_124_256 ();
 FILLCELL_X32 FILLCELL_124_288 ();
 FILLCELL_X32 FILLCELL_124_320 ();
 FILLCELL_X8 FILLCELL_124_352 ();
 FILLCELL_X4 FILLCELL_124_360 ();
 FILLCELL_X32 FILLCELL_124_366 ();
 FILLCELL_X32 FILLCELL_124_398 ();
 FILLCELL_X32 FILLCELL_124_430 ();
 FILLCELL_X32 FILLCELL_124_462 ();
 FILLCELL_X32 FILLCELL_124_494 ();
 FILLCELL_X32 FILLCELL_124_526 ();
 FILLCELL_X32 FILLCELL_124_558 ();
 FILLCELL_X32 FILLCELL_124_590 ();
 FILLCELL_X32 FILLCELL_124_622 ();
 FILLCELL_X32 FILLCELL_124_654 ();
 FILLCELL_X32 FILLCELL_124_686 ();
 FILLCELL_X32 FILLCELL_124_718 ();
 FILLCELL_X32 FILLCELL_124_750 ();
 FILLCELL_X32 FILLCELL_124_782 ();
 FILLCELL_X32 FILLCELL_124_814 ();
 FILLCELL_X32 FILLCELL_124_846 ();
 FILLCELL_X16 FILLCELL_124_878 ();
 FILLCELL_X1 FILLCELL_124_894 ();
 FILLCELL_X32 FILLCELL_124_899 ();
 FILLCELL_X32 FILLCELL_124_931 ();
 FILLCELL_X32 FILLCELL_124_963 ();
 FILLCELL_X32 FILLCELL_124_995 ();
 FILLCELL_X32 FILLCELL_124_1027 ();
 FILLCELL_X32 FILLCELL_124_1059 ();
 FILLCELL_X32 FILLCELL_124_1091 ();
 FILLCELL_X32 FILLCELL_124_1123 ();
 FILLCELL_X32 FILLCELL_124_1155 ();
 FILLCELL_X32 FILLCELL_124_1187 ();
 FILLCELL_X32 FILLCELL_124_1219 ();
 FILLCELL_X32 FILLCELL_124_1251 ();
 FILLCELL_X32 FILLCELL_124_1283 ();
 FILLCELL_X32 FILLCELL_124_1315 ();
 FILLCELL_X32 FILLCELL_124_1347 ();
 FILLCELL_X32 FILLCELL_124_1379 ();
 FILLCELL_X32 FILLCELL_124_1411 ();
 FILLCELL_X32 FILLCELL_124_1443 ();
 FILLCELL_X32 FILLCELL_124_1475 ();
 FILLCELL_X32 FILLCELL_124_1507 ();
 FILLCELL_X32 FILLCELL_124_1539 ();
 FILLCELL_X32 FILLCELL_124_1571 ();
 FILLCELL_X32 FILLCELL_124_1603 ();
 FILLCELL_X32 FILLCELL_124_1635 ();
 FILLCELL_X32 FILLCELL_124_1667 ();
 FILLCELL_X32 FILLCELL_124_1699 ();
 FILLCELL_X32 FILLCELL_124_1731 ();
 FILLCELL_X32 FILLCELL_124_1763 ();
 FILLCELL_X32 FILLCELL_124_1795 ();
 FILLCELL_X32 FILLCELL_124_1827 ();
 FILLCELL_X32 FILLCELL_124_1859 ();
 FILLCELL_X4 FILLCELL_124_1891 ();
 FILLCELL_X2 FILLCELL_124_1895 ();
 FILLCELL_X32 FILLCELL_125_0 ();
 FILLCELL_X32 FILLCELL_125_32 ();
 FILLCELL_X32 FILLCELL_125_64 ();
 FILLCELL_X32 FILLCELL_125_96 ();
 FILLCELL_X16 FILLCELL_125_128 ();
 FILLCELL_X8 FILLCELL_125_144 ();
 FILLCELL_X4 FILLCELL_125_152 ();
 FILLCELL_X2 FILLCELL_125_156 ();
 FILLCELL_X1 FILLCELL_125_158 ();
 FILLCELL_X4 FILLCELL_125_163 ();
 FILLCELL_X2 FILLCELL_125_167 ();
 FILLCELL_X1 FILLCELL_125_169 ();
 FILLCELL_X32 FILLCELL_125_174 ();
 FILLCELL_X32 FILLCELL_125_206 ();
 FILLCELL_X32 FILLCELL_125_238 ();
 FILLCELL_X32 FILLCELL_125_270 ();
 FILLCELL_X32 FILLCELL_125_302 ();
 FILLCELL_X16 FILLCELL_125_334 ();
 FILLCELL_X4 FILLCELL_125_350 ();
 FILLCELL_X2 FILLCELL_125_354 ();
 FILLCELL_X1 FILLCELL_125_356 ();
 FILLCELL_X32 FILLCELL_125_360 ();
 FILLCELL_X32 FILLCELL_125_392 ();
 FILLCELL_X32 FILLCELL_125_424 ();
 FILLCELL_X32 FILLCELL_125_456 ();
 FILLCELL_X32 FILLCELL_125_488 ();
 FILLCELL_X32 FILLCELL_125_520 ();
 FILLCELL_X32 FILLCELL_125_552 ();
 FILLCELL_X32 FILLCELL_125_584 ();
 FILLCELL_X32 FILLCELL_125_616 ();
 FILLCELL_X32 FILLCELL_125_648 ();
 FILLCELL_X32 FILLCELL_125_680 ();
 FILLCELL_X32 FILLCELL_125_712 ();
 FILLCELL_X32 FILLCELL_125_744 ();
 FILLCELL_X32 FILLCELL_125_776 ();
 FILLCELL_X32 FILLCELL_125_808 ();
 FILLCELL_X32 FILLCELL_125_840 ();
 FILLCELL_X32 FILLCELL_125_872 ();
 FILLCELL_X32 FILLCELL_125_904 ();
 FILLCELL_X32 FILLCELL_125_936 ();
 FILLCELL_X32 FILLCELL_125_968 ();
 FILLCELL_X32 FILLCELL_125_1000 ();
 FILLCELL_X32 FILLCELL_125_1032 ();
 FILLCELL_X32 FILLCELL_125_1064 ();
 FILLCELL_X32 FILLCELL_125_1096 ();
 FILLCELL_X32 FILLCELL_125_1128 ();
 FILLCELL_X32 FILLCELL_125_1160 ();
 FILLCELL_X32 FILLCELL_125_1192 ();
 FILLCELL_X32 FILLCELL_125_1224 ();
 FILLCELL_X32 FILLCELL_125_1256 ();
 FILLCELL_X32 FILLCELL_125_1288 ();
 FILLCELL_X32 FILLCELL_125_1320 ();
 FILLCELL_X32 FILLCELL_125_1352 ();
 FILLCELL_X32 FILLCELL_125_1384 ();
 FILLCELL_X32 FILLCELL_125_1416 ();
 FILLCELL_X32 FILLCELL_125_1448 ();
 FILLCELL_X32 FILLCELL_125_1480 ();
 FILLCELL_X32 FILLCELL_125_1512 ();
 FILLCELL_X32 FILLCELL_125_1544 ();
 FILLCELL_X32 FILLCELL_125_1576 ();
 FILLCELL_X32 FILLCELL_125_1608 ();
 FILLCELL_X32 FILLCELL_125_1640 ();
 FILLCELL_X32 FILLCELL_125_1672 ();
 FILLCELL_X32 FILLCELL_125_1704 ();
 FILLCELL_X32 FILLCELL_125_1736 ();
 FILLCELL_X32 FILLCELL_125_1768 ();
 FILLCELL_X32 FILLCELL_125_1800 ();
 FILLCELL_X32 FILLCELL_125_1832 ();
 FILLCELL_X32 FILLCELL_125_1864 ();
 FILLCELL_X1 FILLCELL_125_1896 ();
 FILLCELL_X32 FILLCELL_126_0 ();
 FILLCELL_X32 FILLCELL_126_32 ();
 FILLCELL_X32 FILLCELL_126_64 ();
 FILLCELL_X32 FILLCELL_126_96 ();
 FILLCELL_X32 FILLCELL_126_128 ();
 FILLCELL_X32 FILLCELL_126_160 ();
 FILLCELL_X32 FILLCELL_126_192 ();
 FILLCELL_X4 FILLCELL_126_224 ();
 FILLCELL_X32 FILLCELL_126_231 ();
 FILLCELL_X32 FILLCELL_126_263 ();
 FILLCELL_X32 FILLCELL_126_295 ();
 FILLCELL_X32 FILLCELL_126_327 ();
 FILLCELL_X32 FILLCELL_126_359 ();
 FILLCELL_X32 FILLCELL_126_391 ();
 FILLCELL_X32 FILLCELL_126_423 ();
 FILLCELL_X1 FILLCELL_126_455 ();
 FILLCELL_X32 FILLCELL_126_461 ();
 FILLCELL_X32 FILLCELL_126_493 ();
 FILLCELL_X32 FILLCELL_126_525 ();
 FILLCELL_X8 FILLCELL_126_557 ();
 FILLCELL_X4 FILLCELL_126_565 ();
 FILLCELL_X2 FILLCELL_126_569 ();
 FILLCELL_X32 FILLCELL_126_577 ();
 FILLCELL_X32 FILLCELL_126_609 ();
 FILLCELL_X32 FILLCELL_126_641 ();
 FILLCELL_X32 FILLCELL_126_673 ();
 FILLCELL_X32 FILLCELL_126_705 ();
 FILLCELL_X32 FILLCELL_126_737 ();
 FILLCELL_X32 FILLCELL_126_769 ();
 FILLCELL_X32 FILLCELL_126_801 ();
 FILLCELL_X32 FILLCELL_126_833 ();
 FILLCELL_X32 FILLCELL_126_865 ();
 FILLCELL_X32 FILLCELL_126_897 ();
 FILLCELL_X32 FILLCELL_126_929 ();
 FILLCELL_X32 FILLCELL_126_961 ();
 FILLCELL_X32 FILLCELL_126_993 ();
 FILLCELL_X32 FILLCELL_126_1025 ();
 FILLCELL_X32 FILLCELL_126_1057 ();
 FILLCELL_X32 FILLCELL_126_1089 ();
 FILLCELL_X32 FILLCELL_126_1121 ();
 FILLCELL_X32 FILLCELL_126_1153 ();
 FILLCELL_X32 FILLCELL_126_1185 ();
 FILLCELL_X32 FILLCELL_126_1217 ();
 FILLCELL_X32 FILLCELL_126_1249 ();
 FILLCELL_X32 FILLCELL_126_1281 ();
 FILLCELL_X32 FILLCELL_126_1313 ();
 FILLCELL_X32 FILLCELL_126_1345 ();
 FILLCELL_X32 FILLCELL_126_1377 ();
 FILLCELL_X32 FILLCELL_126_1409 ();
 FILLCELL_X32 FILLCELL_126_1441 ();
 FILLCELL_X32 FILLCELL_126_1473 ();
 FILLCELL_X32 FILLCELL_126_1505 ();
 FILLCELL_X32 FILLCELL_126_1537 ();
 FILLCELL_X32 FILLCELL_126_1569 ();
 FILLCELL_X32 FILLCELL_126_1601 ();
 FILLCELL_X32 FILLCELL_126_1633 ();
 FILLCELL_X32 FILLCELL_126_1665 ();
 FILLCELL_X32 FILLCELL_126_1697 ();
 FILLCELL_X32 FILLCELL_126_1729 ();
 FILLCELL_X32 FILLCELL_126_1761 ();
 FILLCELL_X32 FILLCELL_126_1793 ();
 FILLCELL_X32 FILLCELL_126_1825 ();
 FILLCELL_X32 FILLCELL_126_1857 ();
 FILLCELL_X8 FILLCELL_126_1889 ();
 FILLCELL_X32 FILLCELL_127_0 ();
 FILLCELL_X32 FILLCELL_127_32 ();
 FILLCELL_X32 FILLCELL_127_64 ();
 FILLCELL_X32 FILLCELL_127_96 ();
 FILLCELL_X32 FILLCELL_127_128 ();
 FILLCELL_X32 FILLCELL_127_160 ();
 FILLCELL_X32 FILLCELL_127_192 ();
 FILLCELL_X32 FILLCELL_127_224 ();
 FILLCELL_X32 FILLCELL_127_256 ();
 FILLCELL_X32 FILLCELL_127_288 ();
 FILLCELL_X32 FILLCELL_127_320 ();
 FILLCELL_X32 FILLCELL_127_352 ();
 FILLCELL_X32 FILLCELL_127_384 ();
 FILLCELL_X32 FILLCELL_127_416 ();
 FILLCELL_X32 FILLCELL_127_448 ();
 FILLCELL_X32 FILLCELL_127_480 ();
 FILLCELL_X32 FILLCELL_127_512 ();
 FILLCELL_X2 FILLCELL_127_544 ();
 FILLCELL_X32 FILLCELL_127_548 ();
 FILLCELL_X32 FILLCELL_127_580 ();
 FILLCELL_X4 FILLCELL_127_612 ();
 FILLCELL_X32 FILLCELL_127_620 ();
 FILLCELL_X2 FILLCELL_127_652 ();
 FILLCELL_X32 FILLCELL_127_656 ();
 FILLCELL_X32 FILLCELL_127_688 ();
 FILLCELL_X32 FILLCELL_127_720 ();
 FILLCELL_X32 FILLCELL_127_752 ();
 FILLCELL_X32 FILLCELL_127_784 ();
 FILLCELL_X32 FILLCELL_127_816 ();
 FILLCELL_X32 FILLCELL_127_848 ();
 FILLCELL_X32 FILLCELL_127_880 ();
 FILLCELL_X32 FILLCELL_127_912 ();
 FILLCELL_X32 FILLCELL_127_947 ();
 FILLCELL_X32 FILLCELL_127_979 ();
 FILLCELL_X32 FILLCELL_127_1011 ();
 FILLCELL_X32 FILLCELL_127_1043 ();
 FILLCELL_X32 FILLCELL_127_1075 ();
 FILLCELL_X32 FILLCELL_127_1107 ();
 FILLCELL_X32 FILLCELL_127_1139 ();
 FILLCELL_X32 FILLCELL_127_1171 ();
 FILLCELL_X32 FILLCELL_127_1203 ();
 FILLCELL_X32 FILLCELL_127_1235 ();
 FILLCELL_X32 FILLCELL_127_1267 ();
 FILLCELL_X32 FILLCELL_127_1299 ();
 FILLCELL_X32 FILLCELL_127_1331 ();
 FILLCELL_X32 FILLCELL_127_1363 ();
 FILLCELL_X32 FILLCELL_127_1395 ();
 FILLCELL_X32 FILLCELL_127_1427 ();
 FILLCELL_X32 FILLCELL_127_1459 ();
 FILLCELL_X32 FILLCELL_127_1491 ();
 FILLCELL_X32 FILLCELL_127_1523 ();
 FILLCELL_X32 FILLCELL_127_1555 ();
 FILLCELL_X32 FILLCELL_127_1587 ();
 FILLCELL_X32 FILLCELL_127_1619 ();
 FILLCELL_X32 FILLCELL_127_1651 ();
 FILLCELL_X32 FILLCELL_127_1683 ();
 FILLCELL_X32 FILLCELL_127_1715 ();
 FILLCELL_X32 FILLCELL_127_1747 ();
 FILLCELL_X32 FILLCELL_127_1779 ();
 FILLCELL_X32 FILLCELL_127_1811 ();
 FILLCELL_X32 FILLCELL_127_1843 ();
 FILLCELL_X16 FILLCELL_127_1875 ();
 FILLCELL_X4 FILLCELL_127_1891 ();
 FILLCELL_X2 FILLCELL_127_1895 ();
 FILLCELL_X32 FILLCELL_128_0 ();
 FILLCELL_X32 FILLCELL_128_32 ();
 FILLCELL_X16 FILLCELL_128_64 ();
 FILLCELL_X8 FILLCELL_128_80 ();
 FILLCELL_X2 FILLCELL_128_88 ();
 FILLCELL_X32 FILLCELL_128_92 ();
 FILLCELL_X32 FILLCELL_128_124 ();
 FILLCELL_X32 FILLCELL_128_156 ();
 FILLCELL_X32 FILLCELL_128_188 ();
 FILLCELL_X32 FILLCELL_128_220 ();
 FILLCELL_X4 FILLCELL_128_252 ();
 FILLCELL_X32 FILLCELL_128_260 ();
 FILLCELL_X32 FILLCELL_128_292 ();
 FILLCELL_X32 FILLCELL_128_324 ();
 FILLCELL_X16 FILLCELL_128_356 ();
 FILLCELL_X4 FILLCELL_128_372 ();
 FILLCELL_X2 FILLCELL_128_376 ();
 FILLCELL_X32 FILLCELL_128_381 ();
 FILLCELL_X32 FILLCELL_128_413 ();
 FILLCELL_X32 FILLCELL_128_445 ();
 FILLCELL_X32 FILLCELL_128_477 ();
 FILLCELL_X32 FILLCELL_128_509 ();
 FILLCELL_X32 FILLCELL_128_541 ();
 FILLCELL_X32 FILLCELL_128_573 ();
 FILLCELL_X32 FILLCELL_128_605 ();
 FILLCELL_X32 FILLCELL_128_637 ();
 FILLCELL_X32 FILLCELL_128_669 ();
 FILLCELL_X32 FILLCELL_128_701 ();
 FILLCELL_X32 FILLCELL_128_733 ();
 FILLCELL_X32 FILLCELL_128_765 ();
 FILLCELL_X32 FILLCELL_128_797 ();
 FILLCELL_X32 FILLCELL_128_829 ();
 FILLCELL_X32 FILLCELL_128_861 ();
 FILLCELL_X16 FILLCELL_128_893 ();
 FILLCELL_X32 FILLCELL_128_913 ();
 FILLCELL_X32 FILLCELL_128_945 ();
 FILLCELL_X32 FILLCELL_128_977 ();
 FILLCELL_X32 FILLCELL_128_1009 ();
 FILLCELL_X32 FILLCELL_128_1041 ();
 FILLCELL_X32 FILLCELL_128_1073 ();
 FILLCELL_X32 FILLCELL_128_1105 ();
 FILLCELL_X32 FILLCELL_128_1137 ();
 FILLCELL_X32 FILLCELL_128_1169 ();
 FILLCELL_X32 FILLCELL_128_1201 ();
 FILLCELL_X32 FILLCELL_128_1233 ();
 FILLCELL_X32 FILLCELL_128_1265 ();
 FILLCELL_X32 FILLCELL_128_1297 ();
 FILLCELL_X32 FILLCELL_128_1329 ();
 FILLCELL_X32 FILLCELL_128_1361 ();
 FILLCELL_X32 FILLCELL_128_1393 ();
 FILLCELL_X32 FILLCELL_128_1425 ();
 FILLCELL_X32 FILLCELL_128_1457 ();
 FILLCELL_X32 FILLCELL_128_1489 ();
 FILLCELL_X32 FILLCELL_128_1521 ();
 FILLCELL_X32 FILLCELL_128_1553 ();
 FILLCELL_X32 FILLCELL_128_1585 ();
 FILLCELL_X32 FILLCELL_128_1617 ();
 FILLCELL_X32 FILLCELL_128_1649 ();
 FILLCELL_X32 FILLCELL_128_1681 ();
 FILLCELL_X32 FILLCELL_128_1713 ();
 FILLCELL_X32 FILLCELL_128_1745 ();
 FILLCELL_X32 FILLCELL_128_1777 ();
 FILLCELL_X32 FILLCELL_128_1809 ();
 FILLCELL_X32 FILLCELL_128_1841 ();
 FILLCELL_X16 FILLCELL_128_1873 ();
 FILLCELL_X8 FILLCELL_128_1889 ();
 FILLCELL_X32 FILLCELL_129_0 ();
 FILLCELL_X32 FILLCELL_129_32 ();
 FILLCELL_X32 FILLCELL_129_64 ();
 FILLCELL_X32 FILLCELL_129_96 ();
 FILLCELL_X32 FILLCELL_129_128 ();
 FILLCELL_X32 FILLCELL_129_160 ();
 FILLCELL_X32 FILLCELL_129_192 ();
 FILLCELL_X32 FILLCELL_129_224 ();
 FILLCELL_X32 FILLCELL_129_256 ();
 FILLCELL_X32 FILLCELL_129_288 ();
 FILLCELL_X32 FILLCELL_129_320 ();
 FILLCELL_X16 FILLCELL_129_352 ();
 FILLCELL_X8 FILLCELL_129_368 ();
 FILLCELL_X2 FILLCELL_129_376 ();
 FILLCELL_X1 FILLCELL_129_378 ();
 FILLCELL_X16 FILLCELL_129_382 ();
 FILLCELL_X1 FILLCELL_129_398 ();
 FILLCELL_X32 FILLCELL_129_402 ();
 FILLCELL_X32 FILLCELL_129_434 ();
 FILLCELL_X32 FILLCELL_129_466 ();
 FILLCELL_X32 FILLCELL_129_498 ();
 FILLCELL_X32 FILLCELL_129_530 ();
 FILLCELL_X32 FILLCELL_129_562 ();
 FILLCELL_X32 FILLCELL_129_594 ();
 FILLCELL_X32 FILLCELL_129_626 ();
 FILLCELL_X32 FILLCELL_129_658 ();
 FILLCELL_X32 FILLCELL_129_690 ();
 FILLCELL_X16 FILLCELL_129_722 ();
 FILLCELL_X4 FILLCELL_129_738 ();
 FILLCELL_X2 FILLCELL_129_742 ();
 FILLCELL_X1 FILLCELL_129_744 ();
 FILLCELL_X32 FILLCELL_129_749 ();
 FILLCELL_X32 FILLCELL_129_781 ();
 FILLCELL_X32 FILLCELL_129_813 ();
 FILLCELL_X32 FILLCELL_129_845 ();
 FILLCELL_X32 FILLCELL_129_877 ();
 FILLCELL_X32 FILLCELL_129_909 ();
 FILLCELL_X32 FILLCELL_129_941 ();
 FILLCELL_X32 FILLCELL_129_973 ();
 FILLCELL_X32 FILLCELL_129_1005 ();
 FILLCELL_X32 FILLCELL_129_1037 ();
 FILLCELL_X32 FILLCELL_129_1069 ();
 FILLCELL_X32 FILLCELL_129_1101 ();
 FILLCELL_X32 FILLCELL_129_1133 ();
 FILLCELL_X32 FILLCELL_129_1165 ();
 FILLCELL_X32 FILLCELL_129_1197 ();
 FILLCELL_X32 FILLCELL_129_1229 ();
 FILLCELL_X32 FILLCELL_129_1261 ();
 FILLCELL_X32 FILLCELL_129_1293 ();
 FILLCELL_X32 FILLCELL_129_1325 ();
 FILLCELL_X32 FILLCELL_129_1357 ();
 FILLCELL_X32 FILLCELL_129_1389 ();
 FILLCELL_X32 FILLCELL_129_1421 ();
 FILLCELL_X32 FILLCELL_129_1453 ();
 FILLCELL_X32 FILLCELL_129_1485 ();
 FILLCELL_X32 FILLCELL_129_1517 ();
 FILLCELL_X32 FILLCELL_129_1549 ();
 FILLCELL_X32 FILLCELL_129_1581 ();
 FILLCELL_X32 FILLCELL_129_1613 ();
 FILLCELL_X32 FILLCELL_129_1645 ();
 FILLCELL_X32 FILLCELL_129_1677 ();
 FILLCELL_X32 FILLCELL_129_1709 ();
 FILLCELL_X32 FILLCELL_129_1741 ();
 FILLCELL_X32 FILLCELL_129_1773 ();
 FILLCELL_X32 FILLCELL_129_1805 ();
 FILLCELL_X32 FILLCELL_129_1837 ();
 FILLCELL_X16 FILLCELL_129_1869 ();
 FILLCELL_X8 FILLCELL_129_1885 ();
 FILLCELL_X4 FILLCELL_129_1893 ();
 FILLCELL_X32 FILLCELL_130_0 ();
 FILLCELL_X32 FILLCELL_130_32 ();
 FILLCELL_X32 FILLCELL_130_64 ();
 FILLCELL_X32 FILLCELL_130_96 ();
 FILLCELL_X32 FILLCELL_130_128 ();
 FILLCELL_X32 FILLCELL_130_160 ();
 FILLCELL_X32 FILLCELL_130_192 ();
 FILLCELL_X32 FILLCELL_130_224 ();
 FILLCELL_X32 FILLCELL_130_256 ();
 FILLCELL_X32 FILLCELL_130_288 ();
 FILLCELL_X32 FILLCELL_130_320 ();
 FILLCELL_X32 FILLCELL_130_352 ();
 FILLCELL_X32 FILLCELL_130_384 ();
 FILLCELL_X32 FILLCELL_130_416 ();
 FILLCELL_X32 FILLCELL_130_448 ();
 FILLCELL_X32 FILLCELL_130_480 ();
 FILLCELL_X32 FILLCELL_130_512 ();
 FILLCELL_X32 FILLCELL_130_544 ();
 FILLCELL_X32 FILLCELL_130_576 ();
 FILLCELL_X32 FILLCELL_130_608 ();
 FILLCELL_X32 FILLCELL_130_640 ();
 FILLCELL_X32 FILLCELL_130_672 ();
 FILLCELL_X32 FILLCELL_130_704 ();
 FILLCELL_X32 FILLCELL_130_736 ();
 FILLCELL_X32 FILLCELL_130_768 ();
 FILLCELL_X32 FILLCELL_130_800 ();
 FILLCELL_X32 FILLCELL_130_832 ();
 FILLCELL_X32 FILLCELL_130_864 ();
 FILLCELL_X32 FILLCELL_130_896 ();
 FILLCELL_X32 FILLCELL_130_928 ();
 FILLCELL_X32 FILLCELL_130_960 ();
 FILLCELL_X32 FILLCELL_130_992 ();
 FILLCELL_X32 FILLCELL_130_1024 ();
 FILLCELL_X32 FILLCELL_130_1056 ();
 FILLCELL_X32 FILLCELL_130_1088 ();
 FILLCELL_X8 FILLCELL_130_1120 ();
 FILLCELL_X4 FILLCELL_130_1128 ();
 FILLCELL_X2 FILLCELL_130_1132 ();
 FILLCELL_X1 FILLCELL_130_1134 ();
 FILLCELL_X32 FILLCELL_130_1152 ();
 FILLCELL_X32 FILLCELL_130_1184 ();
 FILLCELL_X32 FILLCELL_130_1216 ();
 FILLCELL_X32 FILLCELL_130_1248 ();
 FILLCELL_X32 FILLCELL_130_1280 ();
 FILLCELL_X32 FILLCELL_130_1312 ();
 FILLCELL_X32 FILLCELL_130_1344 ();
 FILLCELL_X32 FILLCELL_130_1376 ();
 FILLCELL_X32 FILLCELL_130_1408 ();
 FILLCELL_X32 FILLCELL_130_1440 ();
 FILLCELL_X32 FILLCELL_130_1472 ();
 FILLCELL_X32 FILLCELL_130_1504 ();
 FILLCELL_X32 FILLCELL_130_1536 ();
 FILLCELL_X32 FILLCELL_130_1568 ();
 FILLCELL_X32 FILLCELL_130_1600 ();
 FILLCELL_X32 FILLCELL_130_1632 ();
 FILLCELL_X32 FILLCELL_130_1664 ();
 FILLCELL_X32 FILLCELL_130_1696 ();
 FILLCELL_X32 FILLCELL_130_1728 ();
 FILLCELL_X32 FILLCELL_130_1760 ();
 FILLCELL_X32 FILLCELL_130_1792 ();
 FILLCELL_X32 FILLCELL_130_1824 ();
 FILLCELL_X32 FILLCELL_130_1856 ();
 FILLCELL_X8 FILLCELL_130_1888 ();
 FILLCELL_X1 FILLCELL_130_1896 ();
 FILLCELL_X32 FILLCELL_131_0 ();
 FILLCELL_X32 FILLCELL_131_32 ();
 FILLCELL_X32 FILLCELL_131_64 ();
 FILLCELL_X32 FILLCELL_131_96 ();
 FILLCELL_X32 FILLCELL_131_128 ();
 FILLCELL_X32 FILLCELL_131_160 ();
 FILLCELL_X32 FILLCELL_131_192 ();
 FILLCELL_X32 FILLCELL_131_224 ();
 FILLCELL_X32 FILLCELL_131_256 ();
 FILLCELL_X32 FILLCELL_131_292 ();
 FILLCELL_X32 FILLCELL_131_324 ();
 FILLCELL_X32 FILLCELL_131_356 ();
 FILLCELL_X8 FILLCELL_131_388 ();
 FILLCELL_X2 FILLCELL_131_396 ();
 FILLCELL_X32 FILLCELL_131_400 ();
 FILLCELL_X32 FILLCELL_131_432 ();
 FILLCELL_X4 FILLCELL_131_464 ();
 FILLCELL_X2 FILLCELL_131_468 ();
 FILLCELL_X32 FILLCELL_131_472 ();
 FILLCELL_X32 FILLCELL_131_504 ();
 FILLCELL_X32 FILLCELL_131_536 ();
 FILLCELL_X32 FILLCELL_131_573 ();
 FILLCELL_X32 FILLCELL_131_605 ();
 FILLCELL_X32 FILLCELL_131_637 ();
 FILLCELL_X32 FILLCELL_131_669 ();
 FILLCELL_X32 FILLCELL_131_701 ();
 FILLCELL_X16 FILLCELL_131_733 ();
 FILLCELL_X8 FILLCELL_131_749 ();
 FILLCELL_X4 FILLCELL_131_757 ();
 FILLCELL_X2 FILLCELL_131_761 ();
 FILLCELL_X32 FILLCELL_131_767 ();
 FILLCELL_X32 FILLCELL_131_799 ();
 FILLCELL_X32 FILLCELL_131_831 ();
 FILLCELL_X32 FILLCELL_131_863 ();
 FILLCELL_X32 FILLCELL_131_895 ();
 FILLCELL_X32 FILLCELL_131_927 ();
 FILLCELL_X16 FILLCELL_131_959 ();
 FILLCELL_X8 FILLCELL_131_975 ();
 FILLCELL_X2 FILLCELL_131_983 ();
 FILLCELL_X1 FILLCELL_131_985 ();
 FILLCELL_X32 FILLCELL_131_1003 ();
 FILLCELL_X32 FILLCELL_131_1035 ();
 FILLCELL_X16 FILLCELL_131_1067 ();
 FILLCELL_X4 FILLCELL_131_1083 ();
 FILLCELL_X2 FILLCELL_131_1087 ();
 FILLCELL_X1 FILLCELL_131_1089 ();
 FILLCELL_X32 FILLCELL_131_1093 ();
 FILLCELL_X32 FILLCELL_131_1125 ();
 FILLCELL_X32 FILLCELL_131_1157 ();
 FILLCELL_X32 FILLCELL_131_1189 ();
 FILLCELL_X32 FILLCELL_131_1221 ();
 FILLCELL_X32 FILLCELL_131_1253 ();
 FILLCELL_X32 FILLCELL_131_1285 ();
 FILLCELL_X32 FILLCELL_131_1317 ();
 FILLCELL_X32 FILLCELL_131_1349 ();
 FILLCELL_X32 FILLCELL_131_1381 ();
 FILLCELL_X32 FILLCELL_131_1413 ();
 FILLCELL_X32 FILLCELL_131_1445 ();
 FILLCELL_X32 FILLCELL_131_1477 ();
 FILLCELL_X32 FILLCELL_131_1509 ();
 FILLCELL_X32 FILLCELL_131_1541 ();
 FILLCELL_X32 FILLCELL_131_1573 ();
 FILLCELL_X32 FILLCELL_131_1605 ();
 FILLCELL_X32 FILLCELL_131_1637 ();
 FILLCELL_X32 FILLCELL_131_1669 ();
 FILLCELL_X32 FILLCELL_131_1701 ();
 FILLCELL_X32 FILLCELL_131_1733 ();
 FILLCELL_X32 FILLCELL_131_1765 ();
 FILLCELL_X32 FILLCELL_131_1797 ();
 FILLCELL_X32 FILLCELL_131_1829 ();
 FILLCELL_X32 FILLCELL_131_1861 ();
 FILLCELL_X4 FILLCELL_131_1893 ();
 FILLCELL_X32 FILLCELL_132_0 ();
 FILLCELL_X8 FILLCELL_132_32 ();
 FILLCELL_X2 FILLCELL_132_40 ();
 FILLCELL_X32 FILLCELL_132_59 ();
 FILLCELL_X32 FILLCELL_132_91 ();
 FILLCELL_X32 FILLCELL_132_123 ();
 FILLCELL_X32 FILLCELL_132_155 ();
 FILLCELL_X32 FILLCELL_132_187 ();
 FILLCELL_X32 FILLCELL_132_219 ();
 FILLCELL_X32 FILLCELL_132_251 ();
 FILLCELL_X32 FILLCELL_132_283 ();
 FILLCELL_X32 FILLCELL_132_315 ();
 FILLCELL_X32 FILLCELL_132_347 ();
 FILLCELL_X32 FILLCELL_132_379 ();
 FILLCELL_X32 FILLCELL_132_411 ();
 FILLCELL_X8 FILLCELL_132_443 ();
 FILLCELL_X4 FILLCELL_132_451 ();
 FILLCELL_X32 FILLCELL_132_457 ();
 FILLCELL_X32 FILLCELL_132_489 ();
 FILLCELL_X32 FILLCELL_132_521 ();
 FILLCELL_X8 FILLCELL_132_553 ();
 FILLCELL_X1 FILLCELL_132_561 ();
 FILLCELL_X16 FILLCELL_132_570 ();
 FILLCELL_X2 FILLCELL_132_586 ();
 FILLCELL_X32 FILLCELL_132_590 ();
 FILLCELL_X32 FILLCELL_132_622 ();
 FILLCELL_X16 FILLCELL_132_654 ();
 FILLCELL_X4 FILLCELL_132_670 ();
 FILLCELL_X32 FILLCELL_132_678 ();
 FILLCELL_X8 FILLCELL_132_710 ();
 FILLCELL_X2 FILLCELL_132_718 ();
 FILLCELL_X1 FILLCELL_132_720 ();
 FILLCELL_X32 FILLCELL_132_724 ();
 FILLCELL_X4 FILLCELL_132_756 ();
 FILLCELL_X32 FILLCELL_132_769 ();
 FILLCELL_X32 FILLCELL_132_801 ();
 FILLCELL_X32 FILLCELL_132_833 ();
 FILLCELL_X32 FILLCELL_132_865 ();
 FILLCELL_X32 FILLCELL_132_897 ();
 FILLCELL_X32 FILLCELL_132_929 ();
 FILLCELL_X32 FILLCELL_132_961 ();
 FILLCELL_X32 FILLCELL_132_993 ();
 FILLCELL_X32 FILLCELL_132_1025 ();
 FILLCELL_X32 FILLCELL_132_1057 ();
 FILLCELL_X16 FILLCELL_132_1089 ();
 FILLCELL_X32 FILLCELL_132_1112 ();
 FILLCELL_X32 FILLCELL_132_1144 ();
 FILLCELL_X32 FILLCELL_132_1176 ();
 FILLCELL_X32 FILLCELL_132_1208 ();
 FILLCELL_X32 FILLCELL_132_1240 ();
 FILLCELL_X32 FILLCELL_132_1272 ();
 FILLCELL_X32 FILLCELL_132_1304 ();
 FILLCELL_X32 FILLCELL_132_1336 ();
 FILLCELL_X32 FILLCELL_132_1368 ();
 FILLCELL_X32 FILLCELL_132_1400 ();
 FILLCELL_X32 FILLCELL_132_1432 ();
 FILLCELL_X32 FILLCELL_132_1464 ();
 FILLCELL_X32 FILLCELL_132_1496 ();
 FILLCELL_X32 FILLCELL_132_1528 ();
 FILLCELL_X32 FILLCELL_132_1560 ();
 FILLCELL_X32 FILLCELL_132_1592 ();
 FILLCELL_X32 FILLCELL_132_1624 ();
 FILLCELL_X32 FILLCELL_132_1656 ();
 FILLCELL_X32 FILLCELL_132_1688 ();
 FILLCELL_X32 FILLCELL_132_1720 ();
 FILLCELL_X32 FILLCELL_132_1752 ();
 FILLCELL_X32 FILLCELL_132_1784 ();
 FILLCELL_X32 FILLCELL_132_1816 ();
 FILLCELL_X32 FILLCELL_132_1848 ();
 FILLCELL_X16 FILLCELL_132_1880 ();
 FILLCELL_X1 FILLCELL_132_1896 ();
 FILLCELL_X32 FILLCELL_133_0 ();
 FILLCELL_X32 FILLCELL_133_32 ();
 FILLCELL_X32 FILLCELL_133_64 ();
 FILLCELL_X4 FILLCELL_133_96 ();
 FILLCELL_X32 FILLCELL_133_108 ();
 FILLCELL_X32 FILLCELL_133_140 ();
 FILLCELL_X32 FILLCELL_133_172 ();
 FILLCELL_X32 FILLCELL_133_204 ();
 FILLCELL_X32 FILLCELL_133_236 ();
 FILLCELL_X32 FILLCELL_133_268 ();
 FILLCELL_X32 FILLCELL_133_300 ();
 FILLCELL_X32 FILLCELL_133_332 ();
 FILLCELL_X32 FILLCELL_133_364 ();
 FILLCELL_X32 FILLCELL_133_396 ();
 FILLCELL_X32 FILLCELL_133_428 ();
 FILLCELL_X32 FILLCELL_133_460 ();
 FILLCELL_X32 FILLCELL_133_492 ();
 FILLCELL_X32 FILLCELL_133_524 ();
 FILLCELL_X32 FILLCELL_133_556 ();
 FILLCELL_X32 FILLCELL_133_588 ();
 FILLCELL_X32 FILLCELL_133_620 ();
 FILLCELL_X32 FILLCELL_133_652 ();
 FILLCELL_X32 FILLCELL_133_684 ();
 FILLCELL_X32 FILLCELL_133_716 ();
 FILLCELL_X4 FILLCELL_133_748 ();
 FILLCELL_X32 FILLCELL_133_755 ();
 FILLCELL_X32 FILLCELL_133_787 ();
 FILLCELL_X32 FILLCELL_133_819 ();
 FILLCELL_X8 FILLCELL_133_851 ();
 FILLCELL_X4 FILLCELL_133_859 ();
 FILLCELL_X32 FILLCELL_133_868 ();
 FILLCELL_X32 FILLCELL_133_900 ();
 FILLCELL_X32 FILLCELL_133_932 ();
 FILLCELL_X32 FILLCELL_133_964 ();
 FILLCELL_X32 FILLCELL_133_996 ();
 FILLCELL_X32 FILLCELL_133_1028 ();
 FILLCELL_X32 FILLCELL_133_1060 ();
 FILLCELL_X32 FILLCELL_133_1092 ();
 FILLCELL_X32 FILLCELL_133_1124 ();
 FILLCELL_X32 FILLCELL_133_1156 ();
 FILLCELL_X32 FILLCELL_133_1188 ();
 FILLCELL_X32 FILLCELL_133_1220 ();
 FILLCELL_X32 FILLCELL_133_1252 ();
 FILLCELL_X32 FILLCELL_133_1284 ();
 FILLCELL_X32 FILLCELL_133_1316 ();
 FILLCELL_X32 FILLCELL_133_1348 ();
 FILLCELL_X32 FILLCELL_133_1380 ();
 FILLCELL_X32 FILLCELL_133_1412 ();
 FILLCELL_X32 FILLCELL_133_1444 ();
 FILLCELL_X32 FILLCELL_133_1476 ();
 FILLCELL_X32 FILLCELL_133_1508 ();
 FILLCELL_X32 FILLCELL_133_1540 ();
 FILLCELL_X32 FILLCELL_133_1572 ();
 FILLCELL_X32 FILLCELL_133_1604 ();
 FILLCELL_X32 FILLCELL_133_1636 ();
 FILLCELL_X32 FILLCELL_133_1668 ();
 FILLCELL_X32 FILLCELL_133_1700 ();
 FILLCELL_X32 FILLCELL_133_1732 ();
 FILLCELL_X32 FILLCELL_133_1764 ();
 FILLCELL_X32 FILLCELL_133_1796 ();
 FILLCELL_X32 FILLCELL_133_1828 ();
 FILLCELL_X32 FILLCELL_133_1860 ();
 FILLCELL_X4 FILLCELL_133_1892 ();
 FILLCELL_X1 FILLCELL_133_1896 ();
 FILLCELL_X32 FILLCELL_134_0 ();
 FILLCELL_X32 FILLCELL_134_32 ();
 FILLCELL_X32 FILLCELL_134_64 ();
 FILLCELL_X32 FILLCELL_134_96 ();
 FILLCELL_X32 FILLCELL_134_128 ();
 FILLCELL_X32 FILLCELL_134_160 ();
 FILLCELL_X32 FILLCELL_134_192 ();
 FILLCELL_X32 FILLCELL_134_224 ();
 FILLCELL_X32 FILLCELL_134_256 ();
 FILLCELL_X32 FILLCELL_134_288 ();
 FILLCELL_X32 FILLCELL_134_320 ();
 FILLCELL_X32 FILLCELL_134_352 ();
 FILLCELL_X32 FILLCELL_134_384 ();
 FILLCELL_X32 FILLCELL_134_416 ();
 FILLCELL_X32 FILLCELL_134_448 ();
 FILLCELL_X32 FILLCELL_134_480 ();
 FILLCELL_X32 FILLCELL_134_512 ();
 FILLCELL_X32 FILLCELL_134_544 ();
 FILLCELL_X32 FILLCELL_134_576 ();
 FILLCELL_X32 FILLCELL_134_608 ();
 FILLCELL_X32 FILLCELL_134_640 ();
 FILLCELL_X32 FILLCELL_134_672 ();
 FILLCELL_X32 FILLCELL_134_704 ();
 FILLCELL_X32 FILLCELL_134_736 ();
 FILLCELL_X32 FILLCELL_134_768 ();
 FILLCELL_X32 FILLCELL_134_800 ();
 FILLCELL_X32 FILLCELL_134_832 ();
 FILLCELL_X32 FILLCELL_134_864 ();
 FILLCELL_X32 FILLCELL_134_896 ();
 FILLCELL_X32 FILLCELL_134_928 ();
 FILLCELL_X32 FILLCELL_134_960 ();
 FILLCELL_X16 FILLCELL_134_992 ();
 FILLCELL_X4 FILLCELL_134_1008 ();
 FILLCELL_X2 FILLCELL_134_1012 ();
 FILLCELL_X1 FILLCELL_134_1014 ();
 FILLCELL_X32 FILLCELL_134_1017 ();
 FILLCELL_X32 FILLCELL_134_1049 ();
 FILLCELL_X32 FILLCELL_134_1081 ();
 FILLCELL_X32 FILLCELL_134_1113 ();
 FILLCELL_X32 FILLCELL_134_1145 ();
 FILLCELL_X32 FILLCELL_134_1177 ();
 FILLCELL_X32 FILLCELL_134_1209 ();
 FILLCELL_X32 FILLCELL_134_1241 ();
 FILLCELL_X32 FILLCELL_134_1273 ();
 FILLCELL_X32 FILLCELL_134_1305 ();
 FILLCELL_X32 FILLCELL_134_1337 ();
 FILLCELL_X32 FILLCELL_134_1369 ();
 FILLCELL_X32 FILLCELL_134_1401 ();
 FILLCELL_X32 FILLCELL_134_1433 ();
 FILLCELL_X32 FILLCELL_134_1465 ();
 FILLCELL_X32 FILLCELL_134_1497 ();
 FILLCELL_X32 FILLCELL_134_1529 ();
 FILLCELL_X32 FILLCELL_134_1561 ();
 FILLCELL_X32 FILLCELL_134_1593 ();
 FILLCELL_X32 FILLCELL_134_1625 ();
 FILLCELL_X32 FILLCELL_134_1657 ();
 FILLCELL_X32 FILLCELL_134_1689 ();
 FILLCELL_X32 FILLCELL_134_1721 ();
 FILLCELL_X32 FILLCELL_134_1753 ();
 FILLCELL_X32 FILLCELL_134_1785 ();
 FILLCELL_X32 FILLCELL_134_1817 ();
 FILLCELL_X32 FILLCELL_134_1849 ();
 FILLCELL_X16 FILLCELL_134_1881 ();
 FILLCELL_X32 FILLCELL_135_0 ();
 FILLCELL_X32 FILLCELL_135_32 ();
 FILLCELL_X32 FILLCELL_135_64 ();
 FILLCELL_X32 FILLCELL_135_96 ();
 FILLCELL_X16 FILLCELL_135_128 ();
 FILLCELL_X2 FILLCELL_135_144 ();
 FILLCELL_X32 FILLCELL_135_149 ();
 FILLCELL_X32 FILLCELL_135_181 ();
 FILLCELL_X32 FILLCELL_135_213 ();
 FILLCELL_X32 FILLCELL_135_245 ();
 FILLCELL_X32 FILLCELL_135_277 ();
 FILLCELL_X32 FILLCELL_135_309 ();
 FILLCELL_X32 FILLCELL_135_341 ();
 FILLCELL_X32 FILLCELL_135_373 ();
 FILLCELL_X32 FILLCELL_135_405 ();
 FILLCELL_X32 FILLCELL_135_437 ();
 FILLCELL_X32 FILLCELL_135_469 ();
 FILLCELL_X32 FILLCELL_135_501 ();
 FILLCELL_X32 FILLCELL_135_533 ();
 FILLCELL_X32 FILLCELL_135_565 ();
 FILLCELL_X32 FILLCELL_135_597 ();
 FILLCELL_X32 FILLCELL_135_629 ();
 FILLCELL_X32 FILLCELL_135_661 ();
 FILLCELL_X32 FILLCELL_135_693 ();
 FILLCELL_X32 FILLCELL_135_725 ();
 FILLCELL_X32 FILLCELL_135_757 ();
 FILLCELL_X32 FILLCELL_135_789 ();
 FILLCELL_X32 FILLCELL_135_821 ();
 FILLCELL_X8 FILLCELL_135_853 ();
 FILLCELL_X4 FILLCELL_135_861 ();
 FILLCELL_X2 FILLCELL_135_865 ();
 FILLCELL_X32 FILLCELL_135_870 ();
 FILLCELL_X32 FILLCELL_135_902 ();
 FILLCELL_X32 FILLCELL_135_934 ();
 FILLCELL_X8 FILLCELL_135_966 ();
 FILLCELL_X2 FILLCELL_135_974 ();
 FILLCELL_X32 FILLCELL_135_980 ();
 FILLCELL_X1 FILLCELL_135_1012 ();
 FILLCELL_X32 FILLCELL_135_1018 ();
 FILLCELL_X32 FILLCELL_135_1050 ();
 FILLCELL_X32 FILLCELL_135_1082 ();
 FILLCELL_X32 FILLCELL_135_1114 ();
 FILLCELL_X32 FILLCELL_135_1146 ();
 FILLCELL_X32 FILLCELL_135_1178 ();
 FILLCELL_X32 FILLCELL_135_1210 ();
 FILLCELL_X32 FILLCELL_135_1242 ();
 FILLCELL_X32 FILLCELL_135_1274 ();
 FILLCELL_X32 FILLCELL_135_1306 ();
 FILLCELL_X32 FILLCELL_135_1338 ();
 FILLCELL_X32 FILLCELL_135_1370 ();
 FILLCELL_X32 FILLCELL_135_1402 ();
 FILLCELL_X32 FILLCELL_135_1434 ();
 FILLCELL_X32 FILLCELL_135_1466 ();
 FILLCELL_X32 FILLCELL_135_1498 ();
 FILLCELL_X32 FILLCELL_135_1530 ();
 FILLCELL_X32 FILLCELL_135_1562 ();
 FILLCELL_X32 FILLCELL_135_1594 ();
 FILLCELL_X32 FILLCELL_135_1626 ();
 FILLCELL_X32 FILLCELL_135_1658 ();
 FILLCELL_X32 FILLCELL_135_1690 ();
 FILLCELL_X32 FILLCELL_135_1722 ();
 FILLCELL_X32 FILLCELL_135_1754 ();
 FILLCELL_X32 FILLCELL_135_1786 ();
 FILLCELL_X32 FILLCELL_135_1818 ();
 FILLCELL_X32 FILLCELL_135_1850 ();
 FILLCELL_X8 FILLCELL_135_1882 ();
 FILLCELL_X4 FILLCELL_135_1890 ();
 FILLCELL_X2 FILLCELL_135_1894 ();
 FILLCELL_X1 FILLCELL_135_1896 ();
 FILLCELL_X32 FILLCELL_136_0 ();
 FILLCELL_X32 FILLCELL_136_32 ();
 FILLCELL_X32 FILLCELL_136_64 ();
 FILLCELL_X32 FILLCELL_136_96 ();
 FILLCELL_X32 FILLCELL_136_128 ();
 FILLCELL_X32 FILLCELL_136_160 ();
 FILLCELL_X32 FILLCELL_136_192 ();
 FILLCELL_X32 FILLCELL_136_224 ();
 FILLCELL_X32 FILLCELL_136_256 ();
 FILLCELL_X32 FILLCELL_136_288 ();
 FILLCELL_X16 FILLCELL_136_320 ();
 FILLCELL_X2 FILLCELL_136_336 ();
 FILLCELL_X32 FILLCELL_136_341 ();
 FILLCELL_X32 FILLCELL_136_373 ();
 FILLCELL_X32 FILLCELL_136_405 ();
 FILLCELL_X16 FILLCELL_136_437 ();
 FILLCELL_X8 FILLCELL_136_453 ();
 FILLCELL_X4 FILLCELL_136_461 ();
 FILLCELL_X1 FILLCELL_136_465 ();
 FILLCELL_X32 FILLCELL_136_470 ();
 FILLCELL_X16 FILLCELL_136_502 ();
 FILLCELL_X8 FILLCELL_136_518 ();
 FILLCELL_X4 FILLCELL_136_526 ();
 FILLCELL_X1 FILLCELL_136_530 ();
 FILLCELL_X32 FILLCELL_136_534 ();
 FILLCELL_X32 FILLCELL_136_566 ();
 FILLCELL_X32 FILLCELL_136_598 ();
 FILLCELL_X8 FILLCELL_136_630 ();
 FILLCELL_X2 FILLCELL_136_638 ();
 FILLCELL_X1 FILLCELL_136_640 ();
 FILLCELL_X4 FILLCELL_136_646 ();
 FILLCELL_X16 FILLCELL_136_653 ();
 FILLCELL_X8 FILLCELL_136_669 ();
 FILLCELL_X4 FILLCELL_136_677 ();
 FILLCELL_X2 FILLCELL_136_681 ();
 FILLCELL_X1 FILLCELL_136_683 ();
 FILLCELL_X32 FILLCELL_136_687 ();
 FILLCELL_X32 FILLCELL_136_719 ();
 FILLCELL_X32 FILLCELL_136_751 ();
 FILLCELL_X32 FILLCELL_136_783 ();
 FILLCELL_X32 FILLCELL_136_815 ();
 FILLCELL_X4 FILLCELL_136_847 ();
 FILLCELL_X32 FILLCELL_136_855 ();
 FILLCELL_X32 FILLCELL_136_887 ();
 FILLCELL_X32 FILLCELL_136_919 ();
 FILLCELL_X32 FILLCELL_136_951 ();
 FILLCELL_X32 FILLCELL_136_983 ();
 FILLCELL_X32 FILLCELL_136_1015 ();
 FILLCELL_X32 FILLCELL_136_1047 ();
 FILLCELL_X32 FILLCELL_136_1079 ();
 FILLCELL_X32 FILLCELL_136_1111 ();
 FILLCELL_X32 FILLCELL_136_1143 ();
 FILLCELL_X32 FILLCELL_136_1175 ();
 FILLCELL_X32 FILLCELL_136_1207 ();
 FILLCELL_X32 FILLCELL_136_1239 ();
 FILLCELL_X32 FILLCELL_136_1271 ();
 FILLCELL_X32 FILLCELL_136_1303 ();
 FILLCELL_X32 FILLCELL_136_1335 ();
 FILLCELL_X32 FILLCELL_136_1367 ();
 FILLCELL_X32 FILLCELL_136_1399 ();
 FILLCELL_X32 FILLCELL_136_1431 ();
 FILLCELL_X32 FILLCELL_136_1463 ();
 FILLCELL_X32 FILLCELL_136_1495 ();
 FILLCELL_X32 FILLCELL_136_1527 ();
 FILLCELL_X32 FILLCELL_136_1559 ();
 FILLCELL_X32 FILLCELL_136_1591 ();
 FILLCELL_X32 FILLCELL_136_1623 ();
 FILLCELL_X32 FILLCELL_136_1655 ();
 FILLCELL_X32 FILLCELL_136_1687 ();
 FILLCELL_X32 FILLCELL_136_1719 ();
 FILLCELL_X32 FILLCELL_136_1751 ();
 FILLCELL_X32 FILLCELL_136_1783 ();
 FILLCELL_X32 FILLCELL_136_1815 ();
 FILLCELL_X32 FILLCELL_136_1847 ();
 FILLCELL_X16 FILLCELL_136_1879 ();
 FILLCELL_X2 FILLCELL_136_1895 ();
 FILLCELL_X32 FILLCELL_137_0 ();
 FILLCELL_X32 FILLCELL_137_32 ();
 FILLCELL_X8 FILLCELL_137_64 ();
 FILLCELL_X4 FILLCELL_137_72 ();
 FILLCELL_X2 FILLCELL_137_76 ();
 FILLCELL_X8 FILLCELL_137_82 ();
 FILLCELL_X4 FILLCELL_137_90 ();
 FILLCELL_X2 FILLCELL_137_94 ();
 FILLCELL_X1 FILLCELL_137_96 ();
 FILLCELL_X32 FILLCELL_137_99 ();
 FILLCELL_X32 FILLCELL_137_131 ();
 FILLCELL_X32 FILLCELL_137_163 ();
 FILLCELL_X8 FILLCELL_137_195 ();
 FILLCELL_X4 FILLCELL_137_203 ();
 FILLCELL_X2 FILLCELL_137_207 ();
 FILLCELL_X1 FILLCELL_137_209 ();
 FILLCELL_X32 FILLCELL_137_223 ();
 FILLCELL_X32 FILLCELL_137_255 ();
 FILLCELL_X32 FILLCELL_137_287 ();
 FILLCELL_X32 FILLCELL_137_319 ();
 FILLCELL_X32 FILLCELL_137_351 ();
 FILLCELL_X32 FILLCELL_137_383 ();
 FILLCELL_X32 FILLCELL_137_415 ();
 FILLCELL_X32 FILLCELL_137_447 ();
 FILLCELL_X32 FILLCELL_137_479 ();
 FILLCELL_X32 FILLCELL_137_511 ();
 FILLCELL_X32 FILLCELL_137_543 ();
 FILLCELL_X32 FILLCELL_137_575 ();
 FILLCELL_X4 FILLCELL_137_607 ();
 FILLCELL_X2 FILLCELL_137_611 ();
 FILLCELL_X1 FILLCELL_137_613 ();
 FILLCELL_X32 FILLCELL_137_617 ();
 FILLCELL_X32 FILLCELL_137_649 ();
 FILLCELL_X32 FILLCELL_137_681 ();
 FILLCELL_X32 FILLCELL_137_713 ();
 FILLCELL_X32 FILLCELL_137_745 ();
 FILLCELL_X32 FILLCELL_137_777 ();
 FILLCELL_X32 FILLCELL_137_809 ();
 FILLCELL_X32 FILLCELL_137_841 ();
 FILLCELL_X16 FILLCELL_137_873 ();
 FILLCELL_X8 FILLCELL_137_889 ();
 FILLCELL_X2 FILLCELL_137_897 ();
 FILLCELL_X32 FILLCELL_137_901 ();
 FILLCELL_X32 FILLCELL_137_933 ();
 FILLCELL_X32 FILLCELL_137_965 ();
 FILLCELL_X32 FILLCELL_137_997 ();
 FILLCELL_X32 FILLCELL_137_1029 ();
 FILLCELL_X32 FILLCELL_137_1061 ();
 FILLCELL_X32 FILLCELL_137_1093 ();
 FILLCELL_X32 FILLCELL_137_1125 ();
 FILLCELL_X32 FILLCELL_137_1157 ();
 FILLCELL_X32 FILLCELL_137_1189 ();
 FILLCELL_X32 FILLCELL_137_1221 ();
 FILLCELL_X32 FILLCELL_137_1253 ();
 FILLCELL_X32 FILLCELL_137_1285 ();
 FILLCELL_X32 FILLCELL_137_1317 ();
 FILLCELL_X32 FILLCELL_137_1349 ();
 FILLCELL_X32 FILLCELL_137_1381 ();
 FILLCELL_X32 FILLCELL_137_1413 ();
 FILLCELL_X32 FILLCELL_137_1445 ();
 FILLCELL_X32 FILLCELL_137_1477 ();
 FILLCELL_X32 FILLCELL_137_1509 ();
 FILLCELL_X32 FILLCELL_137_1541 ();
 FILLCELL_X32 FILLCELL_137_1573 ();
 FILLCELL_X32 FILLCELL_137_1605 ();
 FILLCELL_X32 FILLCELL_137_1637 ();
 FILLCELL_X32 FILLCELL_137_1669 ();
 FILLCELL_X32 FILLCELL_137_1701 ();
 FILLCELL_X32 FILLCELL_137_1733 ();
 FILLCELL_X32 FILLCELL_137_1765 ();
 FILLCELL_X32 FILLCELL_137_1797 ();
 FILLCELL_X32 FILLCELL_137_1829 ();
 FILLCELL_X32 FILLCELL_137_1861 ();
 FILLCELL_X4 FILLCELL_137_1893 ();
 FILLCELL_X32 FILLCELL_138_0 ();
 FILLCELL_X32 FILLCELL_138_32 ();
 FILLCELL_X32 FILLCELL_138_64 ();
 FILLCELL_X32 FILLCELL_138_96 ();
 FILLCELL_X32 FILLCELL_138_128 ();
 FILLCELL_X32 FILLCELL_138_160 ();
 FILLCELL_X32 FILLCELL_138_192 ();
 FILLCELL_X32 FILLCELL_138_224 ();
 FILLCELL_X32 FILLCELL_138_256 ();
 FILLCELL_X8 FILLCELL_138_288 ();
 FILLCELL_X2 FILLCELL_138_296 ();
 FILLCELL_X32 FILLCELL_138_311 ();
 FILLCELL_X32 FILLCELL_138_343 ();
 FILLCELL_X32 FILLCELL_138_375 ();
 FILLCELL_X32 FILLCELL_138_407 ();
 FILLCELL_X8 FILLCELL_138_439 ();
 FILLCELL_X2 FILLCELL_138_447 ();
 FILLCELL_X1 FILLCELL_138_449 ();
 FILLCELL_X4 FILLCELL_138_455 ();
 FILLCELL_X1 FILLCELL_138_459 ();
 FILLCELL_X2 FILLCELL_138_464 ();
 FILLCELL_X32 FILLCELL_138_471 ();
 FILLCELL_X32 FILLCELL_138_503 ();
 FILLCELL_X1 FILLCELL_138_535 ();
 FILLCELL_X32 FILLCELL_138_539 ();
 FILLCELL_X32 FILLCELL_138_571 ();
 FILLCELL_X32 FILLCELL_138_603 ();
 FILLCELL_X32 FILLCELL_138_635 ();
 FILLCELL_X32 FILLCELL_138_667 ();
 FILLCELL_X32 FILLCELL_138_699 ();
 FILLCELL_X32 FILLCELL_138_731 ();
 FILLCELL_X32 FILLCELL_138_763 ();
 FILLCELL_X32 FILLCELL_138_795 ();
 FILLCELL_X8 FILLCELL_138_827 ();
 FILLCELL_X4 FILLCELL_138_835 ();
 FILLCELL_X2 FILLCELL_138_839 ();
 FILLCELL_X32 FILLCELL_138_846 ();
 FILLCELL_X8 FILLCELL_138_878 ();
 FILLCELL_X1 FILLCELL_138_886 ();
 FILLCELL_X32 FILLCELL_138_892 ();
 FILLCELL_X32 FILLCELL_138_924 ();
 FILLCELL_X32 FILLCELL_138_956 ();
 FILLCELL_X32 FILLCELL_138_988 ();
 FILLCELL_X32 FILLCELL_138_1020 ();
 FILLCELL_X32 FILLCELL_138_1052 ();
 FILLCELL_X32 FILLCELL_138_1084 ();
 FILLCELL_X32 FILLCELL_138_1116 ();
 FILLCELL_X32 FILLCELL_138_1148 ();
 FILLCELL_X32 FILLCELL_138_1180 ();
 FILLCELL_X32 FILLCELL_138_1212 ();
 FILLCELL_X32 FILLCELL_138_1244 ();
 FILLCELL_X32 FILLCELL_138_1276 ();
 FILLCELL_X32 FILLCELL_138_1308 ();
 FILLCELL_X32 FILLCELL_138_1340 ();
 FILLCELL_X32 FILLCELL_138_1372 ();
 FILLCELL_X32 FILLCELL_138_1404 ();
 FILLCELL_X32 FILLCELL_138_1436 ();
 FILLCELL_X32 FILLCELL_138_1468 ();
 FILLCELL_X32 FILLCELL_138_1500 ();
 FILLCELL_X32 FILLCELL_138_1532 ();
 FILLCELL_X32 FILLCELL_138_1564 ();
 FILLCELL_X32 FILLCELL_138_1596 ();
 FILLCELL_X32 FILLCELL_138_1628 ();
 FILLCELL_X32 FILLCELL_138_1660 ();
 FILLCELL_X32 FILLCELL_138_1692 ();
 FILLCELL_X32 FILLCELL_138_1724 ();
 FILLCELL_X32 FILLCELL_138_1756 ();
 FILLCELL_X32 FILLCELL_138_1788 ();
 FILLCELL_X32 FILLCELL_138_1820 ();
 FILLCELL_X32 FILLCELL_138_1852 ();
 FILLCELL_X8 FILLCELL_138_1884 ();
 FILLCELL_X4 FILLCELL_138_1892 ();
 FILLCELL_X1 FILLCELL_138_1896 ();
 FILLCELL_X32 FILLCELL_139_0 ();
 FILLCELL_X32 FILLCELL_139_32 ();
 FILLCELL_X32 FILLCELL_139_64 ();
 FILLCELL_X32 FILLCELL_139_96 ();
 FILLCELL_X32 FILLCELL_139_128 ();
 FILLCELL_X32 FILLCELL_139_160 ();
 FILLCELL_X32 FILLCELL_139_192 ();
 FILLCELL_X32 FILLCELL_139_224 ();
 FILLCELL_X32 FILLCELL_139_256 ();
 FILLCELL_X32 FILLCELL_139_288 ();
 FILLCELL_X32 FILLCELL_139_320 ();
 FILLCELL_X32 FILLCELL_139_352 ();
 FILLCELL_X32 FILLCELL_139_384 ();
 FILLCELL_X32 FILLCELL_139_416 ();
 FILLCELL_X32 FILLCELL_139_448 ();
 FILLCELL_X32 FILLCELL_139_480 ();
 FILLCELL_X32 FILLCELL_139_512 ();
 FILLCELL_X32 FILLCELL_139_544 ();
 FILLCELL_X32 FILLCELL_139_576 ();
 FILLCELL_X32 FILLCELL_139_608 ();
 FILLCELL_X32 FILLCELL_139_640 ();
 FILLCELL_X32 FILLCELL_139_672 ();
 FILLCELL_X32 FILLCELL_139_704 ();
 FILLCELL_X32 FILLCELL_139_736 ();
 FILLCELL_X32 FILLCELL_139_768 ();
 FILLCELL_X32 FILLCELL_139_800 ();
 FILLCELL_X32 FILLCELL_139_832 ();
 FILLCELL_X32 FILLCELL_139_864 ();
 FILLCELL_X32 FILLCELL_139_896 ();
 FILLCELL_X32 FILLCELL_139_928 ();
 FILLCELL_X32 FILLCELL_139_960 ();
 FILLCELL_X32 FILLCELL_139_992 ();
 FILLCELL_X32 FILLCELL_139_1024 ();
 FILLCELL_X16 FILLCELL_139_1056 ();
 FILLCELL_X8 FILLCELL_139_1072 ();
 FILLCELL_X4 FILLCELL_139_1080 ();
 FILLCELL_X2 FILLCELL_139_1084 ();
 FILLCELL_X8 FILLCELL_139_1090 ();
 FILLCELL_X1 FILLCELL_139_1098 ();
 FILLCELL_X32 FILLCELL_139_1102 ();
 FILLCELL_X32 FILLCELL_139_1134 ();
 FILLCELL_X32 FILLCELL_139_1166 ();
 FILLCELL_X32 FILLCELL_139_1198 ();
 FILLCELL_X32 FILLCELL_139_1230 ();
 FILLCELL_X32 FILLCELL_139_1262 ();
 FILLCELL_X32 FILLCELL_139_1294 ();
 FILLCELL_X32 FILLCELL_139_1326 ();
 FILLCELL_X32 FILLCELL_139_1358 ();
 FILLCELL_X32 FILLCELL_139_1390 ();
 FILLCELL_X32 FILLCELL_139_1422 ();
 FILLCELL_X32 FILLCELL_139_1454 ();
 FILLCELL_X32 FILLCELL_139_1486 ();
 FILLCELL_X32 FILLCELL_139_1518 ();
 FILLCELL_X32 FILLCELL_139_1550 ();
 FILLCELL_X32 FILLCELL_139_1582 ();
 FILLCELL_X32 FILLCELL_139_1614 ();
 FILLCELL_X32 FILLCELL_139_1646 ();
 FILLCELL_X32 FILLCELL_139_1678 ();
 FILLCELL_X32 FILLCELL_139_1710 ();
 FILLCELL_X32 FILLCELL_139_1742 ();
 FILLCELL_X32 FILLCELL_139_1774 ();
 FILLCELL_X32 FILLCELL_139_1806 ();
 FILLCELL_X32 FILLCELL_139_1838 ();
 FILLCELL_X16 FILLCELL_139_1870 ();
 FILLCELL_X8 FILLCELL_139_1886 ();
 FILLCELL_X2 FILLCELL_139_1894 ();
 FILLCELL_X1 FILLCELL_139_1896 ();
 FILLCELL_X32 FILLCELL_140_0 ();
 FILLCELL_X32 FILLCELL_140_32 ();
 FILLCELL_X32 FILLCELL_140_64 ();
 FILLCELL_X32 FILLCELL_140_96 ();
 FILLCELL_X32 FILLCELL_140_128 ();
 FILLCELL_X32 FILLCELL_140_160 ();
 FILLCELL_X16 FILLCELL_140_192 ();
 FILLCELL_X8 FILLCELL_140_208 ();
 FILLCELL_X4 FILLCELL_140_216 ();
 FILLCELL_X32 FILLCELL_140_222 ();
 FILLCELL_X32 FILLCELL_140_254 ();
 FILLCELL_X32 FILLCELL_140_286 ();
 FILLCELL_X32 FILLCELL_140_318 ();
 FILLCELL_X16 FILLCELL_140_350 ();
 FILLCELL_X2 FILLCELL_140_366 ();
 FILLCELL_X1 FILLCELL_140_368 ();
 FILLCELL_X32 FILLCELL_140_378 ();
 FILLCELL_X32 FILLCELL_140_410 ();
 FILLCELL_X32 FILLCELL_140_442 ();
 FILLCELL_X32 FILLCELL_140_474 ();
 FILLCELL_X32 FILLCELL_140_506 ();
 FILLCELL_X32 FILLCELL_140_538 ();
 FILLCELL_X32 FILLCELL_140_570 ();
 FILLCELL_X32 FILLCELL_140_602 ();
 FILLCELL_X4 FILLCELL_140_634 ();
 FILLCELL_X2 FILLCELL_140_638 ();
 FILLCELL_X1 FILLCELL_140_640 ();
 FILLCELL_X32 FILLCELL_140_647 ();
 FILLCELL_X32 FILLCELL_140_679 ();
 FILLCELL_X32 FILLCELL_140_711 ();
 FILLCELL_X32 FILLCELL_140_743 ();
 FILLCELL_X32 FILLCELL_140_775 ();
 FILLCELL_X32 FILLCELL_140_807 ();
 FILLCELL_X16 FILLCELL_140_839 ();
 FILLCELL_X4 FILLCELL_140_855 ();
 FILLCELL_X1 FILLCELL_140_859 ();
 FILLCELL_X16 FILLCELL_140_862 ();
 FILLCELL_X8 FILLCELL_140_878 ();
 FILLCELL_X1 FILLCELL_140_886 ();
 FILLCELL_X32 FILLCELL_140_890 ();
 FILLCELL_X32 FILLCELL_140_922 ();
 FILLCELL_X32 FILLCELL_140_954 ();
 FILLCELL_X32 FILLCELL_140_986 ();
 FILLCELL_X32 FILLCELL_140_1018 ();
 FILLCELL_X32 FILLCELL_140_1050 ();
 FILLCELL_X32 FILLCELL_140_1082 ();
 FILLCELL_X32 FILLCELL_140_1114 ();
 FILLCELL_X32 FILLCELL_140_1146 ();
 FILLCELL_X32 FILLCELL_140_1178 ();
 FILLCELL_X32 FILLCELL_140_1210 ();
 FILLCELL_X32 FILLCELL_140_1242 ();
 FILLCELL_X32 FILLCELL_140_1274 ();
 FILLCELL_X32 FILLCELL_140_1306 ();
 FILLCELL_X32 FILLCELL_140_1338 ();
 FILLCELL_X32 FILLCELL_140_1370 ();
 FILLCELL_X32 FILLCELL_140_1402 ();
 FILLCELL_X32 FILLCELL_140_1434 ();
 FILLCELL_X32 FILLCELL_140_1466 ();
 FILLCELL_X32 FILLCELL_140_1498 ();
 FILLCELL_X32 FILLCELL_140_1530 ();
 FILLCELL_X32 FILLCELL_140_1562 ();
 FILLCELL_X32 FILLCELL_140_1594 ();
 FILLCELL_X32 FILLCELL_140_1626 ();
 FILLCELL_X32 FILLCELL_140_1658 ();
 FILLCELL_X32 FILLCELL_140_1690 ();
 FILLCELL_X32 FILLCELL_140_1722 ();
 FILLCELL_X32 FILLCELL_140_1754 ();
 FILLCELL_X32 FILLCELL_140_1786 ();
 FILLCELL_X32 FILLCELL_140_1818 ();
 FILLCELL_X32 FILLCELL_140_1850 ();
 FILLCELL_X8 FILLCELL_140_1882 ();
 FILLCELL_X4 FILLCELL_140_1890 ();
 FILLCELL_X2 FILLCELL_140_1894 ();
 FILLCELL_X1 FILLCELL_140_1896 ();
 FILLCELL_X32 FILLCELL_141_0 ();
 FILLCELL_X32 FILLCELL_141_32 ();
 FILLCELL_X32 FILLCELL_141_64 ();
 FILLCELL_X32 FILLCELL_141_96 ();
 FILLCELL_X32 FILLCELL_141_128 ();
 FILLCELL_X32 FILLCELL_141_160 ();
 FILLCELL_X32 FILLCELL_141_192 ();
 FILLCELL_X32 FILLCELL_141_224 ();
 FILLCELL_X32 FILLCELL_141_256 ();
 FILLCELL_X32 FILLCELL_141_288 ();
 FILLCELL_X32 FILLCELL_141_320 ();
 FILLCELL_X32 FILLCELL_141_352 ();
 FILLCELL_X32 FILLCELL_141_384 ();
 FILLCELL_X32 FILLCELL_141_416 ();
 FILLCELL_X32 FILLCELL_141_448 ();
 FILLCELL_X32 FILLCELL_141_480 ();
 FILLCELL_X32 FILLCELL_141_512 ();
 FILLCELL_X32 FILLCELL_141_544 ();
 FILLCELL_X32 FILLCELL_141_576 ();
 FILLCELL_X32 FILLCELL_141_608 ();
 FILLCELL_X32 FILLCELL_141_640 ();
 FILLCELL_X32 FILLCELL_141_672 ();
 FILLCELL_X32 FILLCELL_141_704 ();
 FILLCELL_X32 FILLCELL_141_736 ();
 FILLCELL_X32 FILLCELL_141_768 ();
 FILLCELL_X32 FILLCELL_141_800 ();
 FILLCELL_X32 FILLCELL_141_832 ();
 FILLCELL_X32 FILLCELL_141_864 ();
 FILLCELL_X32 FILLCELL_141_896 ();
 FILLCELL_X32 FILLCELL_141_928 ();
 FILLCELL_X32 FILLCELL_141_960 ();
 FILLCELL_X32 FILLCELL_141_992 ();
 FILLCELL_X32 FILLCELL_141_1024 ();
 FILLCELL_X32 FILLCELL_141_1056 ();
 FILLCELL_X32 FILLCELL_141_1088 ();
 FILLCELL_X32 FILLCELL_141_1120 ();
 FILLCELL_X32 FILLCELL_141_1152 ();
 FILLCELL_X32 FILLCELL_141_1184 ();
 FILLCELL_X32 FILLCELL_141_1216 ();
 FILLCELL_X32 FILLCELL_141_1248 ();
 FILLCELL_X32 FILLCELL_141_1280 ();
 FILLCELL_X32 FILLCELL_141_1312 ();
 FILLCELL_X32 FILLCELL_141_1344 ();
 FILLCELL_X32 FILLCELL_141_1376 ();
 FILLCELL_X32 FILLCELL_141_1408 ();
 FILLCELL_X32 FILLCELL_141_1440 ();
 FILLCELL_X32 FILLCELL_141_1472 ();
 FILLCELL_X32 FILLCELL_141_1504 ();
 FILLCELL_X32 FILLCELL_141_1536 ();
 FILLCELL_X32 FILLCELL_141_1568 ();
 FILLCELL_X32 FILLCELL_141_1600 ();
 FILLCELL_X32 FILLCELL_141_1632 ();
 FILLCELL_X32 FILLCELL_141_1664 ();
 FILLCELL_X32 FILLCELL_141_1696 ();
 FILLCELL_X32 FILLCELL_141_1728 ();
 FILLCELL_X32 FILLCELL_141_1760 ();
 FILLCELL_X32 FILLCELL_141_1792 ();
 FILLCELL_X32 FILLCELL_141_1824 ();
 FILLCELL_X32 FILLCELL_141_1856 ();
 FILLCELL_X8 FILLCELL_141_1888 ();
 FILLCELL_X1 FILLCELL_141_1896 ();
 FILLCELL_X32 FILLCELL_142_0 ();
 FILLCELL_X32 FILLCELL_142_32 ();
 FILLCELL_X32 FILLCELL_142_64 ();
 FILLCELL_X32 FILLCELL_142_96 ();
 FILLCELL_X32 FILLCELL_142_128 ();
 FILLCELL_X32 FILLCELL_142_160 ();
 FILLCELL_X32 FILLCELL_142_192 ();
 FILLCELL_X32 FILLCELL_142_224 ();
 FILLCELL_X32 FILLCELL_142_256 ();
 FILLCELL_X32 FILLCELL_142_288 ();
 FILLCELL_X32 FILLCELL_142_320 ();
 FILLCELL_X32 FILLCELL_142_352 ();
 FILLCELL_X32 FILLCELL_142_384 ();
 FILLCELL_X32 FILLCELL_142_416 ();
 FILLCELL_X32 FILLCELL_142_448 ();
 FILLCELL_X32 FILLCELL_142_480 ();
 FILLCELL_X32 FILLCELL_142_512 ();
 FILLCELL_X32 FILLCELL_142_544 ();
 FILLCELL_X32 FILLCELL_142_576 ();
 FILLCELL_X32 FILLCELL_142_608 ();
 FILLCELL_X32 FILLCELL_142_640 ();
 FILLCELL_X32 FILLCELL_142_672 ();
 FILLCELL_X32 FILLCELL_142_704 ();
 FILLCELL_X32 FILLCELL_142_736 ();
 FILLCELL_X16 FILLCELL_142_768 ();
 FILLCELL_X2 FILLCELL_142_784 ();
 FILLCELL_X16 FILLCELL_142_788 ();
 FILLCELL_X1 FILLCELL_142_804 ();
 FILLCELL_X32 FILLCELL_142_807 ();
 FILLCELL_X32 FILLCELL_142_839 ();
 FILLCELL_X4 FILLCELL_142_871 ();
 FILLCELL_X2 FILLCELL_142_875 ();
 FILLCELL_X32 FILLCELL_142_880 ();
 FILLCELL_X32 FILLCELL_142_912 ();
 FILLCELL_X32 FILLCELL_142_944 ();
 FILLCELL_X32 FILLCELL_142_976 ();
 FILLCELL_X32 FILLCELL_142_1008 ();
 FILLCELL_X32 FILLCELL_142_1040 ();
 FILLCELL_X32 FILLCELL_142_1072 ();
 FILLCELL_X32 FILLCELL_142_1104 ();
 FILLCELL_X32 FILLCELL_142_1136 ();
 FILLCELL_X32 FILLCELL_142_1168 ();
 FILLCELL_X32 FILLCELL_142_1200 ();
 FILLCELL_X32 FILLCELL_142_1232 ();
 FILLCELL_X32 FILLCELL_142_1264 ();
 FILLCELL_X32 FILLCELL_142_1296 ();
 FILLCELL_X32 FILLCELL_142_1328 ();
 FILLCELL_X32 FILLCELL_142_1360 ();
 FILLCELL_X32 FILLCELL_142_1392 ();
 FILLCELL_X32 FILLCELL_142_1424 ();
 FILLCELL_X32 FILLCELL_142_1456 ();
 FILLCELL_X32 FILLCELL_142_1488 ();
 FILLCELL_X32 FILLCELL_142_1520 ();
 FILLCELL_X32 FILLCELL_142_1552 ();
 FILLCELL_X32 FILLCELL_142_1584 ();
 FILLCELL_X32 FILLCELL_142_1616 ();
 FILLCELL_X32 FILLCELL_142_1648 ();
 FILLCELL_X32 FILLCELL_142_1680 ();
 FILLCELL_X32 FILLCELL_142_1712 ();
 FILLCELL_X32 FILLCELL_142_1744 ();
 FILLCELL_X32 FILLCELL_142_1776 ();
 FILLCELL_X32 FILLCELL_142_1808 ();
 FILLCELL_X32 FILLCELL_142_1840 ();
 FILLCELL_X16 FILLCELL_142_1872 ();
 FILLCELL_X8 FILLCELL_142_1888 ();
 FILLCELL_X1 FILLCELL_142_1896 ();
 FILLCELL_X32 FILLCELL_143_0 ();
 FILLCELL_X32 FILLCELL_143_32 ();
 FILLCELL_X32 FILLCELL_143_64 ();
 FILLCELL_X32 FILLCELL_143_96 ();
 FILLCELL_X32 FILLCELL_143_128 ();
 FILLCELL_X32 FILLCELL_143_160 ();
 FILLCELL_X32 FILLCELL_143_192 ();
 FILLCELL_X32 FILLCELL_143_224 ();
 FILLCELL_X32 FILLCELL_143_256 ();
 FILLCELL_X32 FILLCELL_143_288 ();
 FILLCELL_X32 FILLCELL_143_320 ();
 FILLCELL_X32 FILLCELL_143_352 ();
 FILLCELL_X32 FILLCELL_143_384 ();
 FILLCELL_X32 FILLCELL_143_416 ();
 FILLCELL_X32 FILLCELL_143_448 ();
 FILLCELL_X32 FILLCELL_143_480 ();
 FILLCELL_X32 FILLCELL_143_512 ();
 FILLCELL_X32 FILLCELL_143_544 ();
 FILLCELL_X32 FILLCELL_143_576 ();
 FILLCELL_X32 FILLCELL_143_608 ();
 FILLCELL_X32 FILLCELL_143_640 ();
 FILLCELL_X32 FILLCELL_143_672 ();
 FILLCELL_X32 FILLCELL_143_704 ();
 FILLCELL_X32 FILLCELL_143_736 ();
 FILLCELL_X32 FILLCELL_143_768 ();
 FILLCELL_X32 FILLCELL_143_800 ();
 FILLCELL_X32 FILLCELL_143_832 ();
 FILLCELL_X32 FILLCELL_143_864 ();
 FILLCELL_X32 FILLCELL_143_896 ();
 FILLCELL_X32 FILLCELL_143_928 ();
 FILLCELL_X32 FILLCELL_143_960 ();
 FILLCELL_X32 FILLCELL_143_992 ();
 FILLCELL_X32 FILLCELL_143_1024 ();
 FILLCELL_X32 FILLCELL_143_1056 ();
 FILLCELL_X16 FILLCELL_143_1088 ();
 FILLCELL_X8 FILLCELL_143_1104 ();
 FILLCELL_X4 FILLCELL_143_1112 ();
 FILLCELL_X32 FILLCELL_143_1119 ();
 FILLCELL_X32 FILLCELL_143_1151 ();
 FILLCELL_X32 FILLCELL_143_1183 ();
 FILLCELL_X32 FILLCELL_143_1215 ();
 FILLCELL_X32 FILLCELL_143_1247 ();
 FILLCELL_X32 FILLCELL_143_1279 ();
 FILLCELL_X32 FILLCELL_143_1311 ();
 FILLCELL_X32 FILLCELL_143_1343 ();
 FILLCELL_X32 FILLCELL_143_1375 ();
 FILLCELL_X32 FILLCELL_143_1407 ();
 FILLCELL_X32 FILLCELL_143_1439 ();
 FILLCELL_X32 FILLCELL_143_1471 ();
 FILLCELL_X32 FILLCELL_143_1503 ();
 FILLCELL_X32 FILLCELL_143_1535 ();
 FILLCELL_X32 FILLCELL_143_1567 ();
 FILLCELL_X32 FILLCELL_143_1599 ();
 FILLCELL_X32 FILLCELL_143_1631 ();
 FILLCELL_X32 FILLCELL_143_1663 ();
 FILLCELL_X32 FILLCELL_143_1695 ();
 FILLCELL_X32 FILLCELL_143_1727 ();
 FILLCELL_X32 FILLCELL_143_1759 ();
 FILLCELL_X32 FILLCELL_143_1791 ();
 FILLCELL_X32 FILLCELL_143_1823 ();
 FILLCELL_X32 FILLCELL_143_1855 ();
 FILLCELL_X8 FILLCELL_143_1887 ();
 FILLCELL_X2 FILLCELL_143_1895 ();
 FILLCELL_X32 FILLCELL_144_0 ();
 FILLCELL_X32 FILLCELL_144_32 ();
 FILLCELL_X16 FILLCELL_144_64 ();
 FILLCELL_X32 FILLCELL_144_84 ();
 FILLCELL_X32 FILLCELL_144_116 ();
 FILLCELL_X32 FILLCELL_144_148 ();
 FILLCELL_X32 FILLCELL_144_180 ();
 FILLCELL_X32 FILLCELL_144_212 ();
 FILLCELL_X32 FILLCELL_144_244 ();
 FILLCELL_X32 FILLCELL_144_276 ();
 FILLCELL_X32 FILLCELL_144_308 ();
 FILLCELL_X32 FILLCELL_144_340 ();
 FILLCELL_X32 FILLCELL_144_372 ();
 FILLCELL_X32 FILLCELL_144_404 ();
 FILLCELL_X32 FILLCELL_144_436 ();
 FILLCELL_X32 FILLCELL_144_468 ();
 FILLCELL_X32 FILLCELL_144_500 ();
 FILLCELL_X32 FILLCELL_144_532 ();
 FILLCELL_X32 FILLCELL_144_564 ();
 FILLCELL_X32 FILLCELL_144_596 ();
 FILLCELL_X32 FILLCELL_144_628 ();
 FILLCELL_X32 FILLCELL_144_660 ();
 FILLCELL_X32 FILLCELL_144_692 ();
 FILLCELL_X32 FILLCELL_144_724 ();
 FILLCELL_X32 FILLCELL_144_756 ();
 FILLCELL_X32 FILLCELL_144_788 ();
 FILLCELL_X32 FILLCELL_144_820 ();
 FILLCELL_X32 FILLCELL_144_852 ();
 FILLCELL_X32 FILLCELL_144_884 ();
 FILLCELL_X32 FILLCELL_144_916 ();
 FILLCELL_X32 FILLCELL_144_948 ();
 FILLCELL_X32 FILLCELL_144_980 ();
 FILLCELL_X32 FILLCELL_144_1012 ();
 FILLCELL_X32 FILLCELL_144_1044 ();
 FILLCELL_X32 FILLCELL_144_1076 ();
 FILLCELL_X8 FILLCELL_144_1108 ();
 FILLCELL_X32 FILLCELL_144_1119 ();
 FILLCELL_X32 FILLCELL_144_1151 ();
 FILLCELL_X32 FILLCELL_144_1183 ();
 FILLCELL_X32 FILLCELL_144_1215 ();
 FILLCELL_X32 FILLCELL_144_1247 ();
 FILLCELL_X32 FILLCELL_144_1279 ();
 FILLCELL_X32 FILLCELL_144_1311 ();
 FILLCELL_X32 FILLCELL_144_1343 ();
 FILLCELL_X32 FILLCELL_144_1375 ();
 FILLCELL_X32 FILLCELL_144_1407 ();
 FILLCELL_X32 FILLCELL_144_1439 ();
 FILLCELL_X32 FILLCELL_144_1471 ();
 FILLCELL_X32 FILLCELL_144_1503 ();
 FILLCELL_X32 FILLCELL_144_1535 ();
 FILLCELL_X32 FILLCELL_144_1567 ();
 FILLCELL_X32 FILLCELL_144_1599 ();
 FILLCELL_X32 FILLCELL_144_1631 ();
 FILLCELL_X32 FILLCELL_144_1663 ();
 FILLCELL_X32 FILLCELL_144_1695 ();
 FILLCELL_X32 FILLCELL_144_1727 ();
 FILLCELL_X32 FILLCELL_144_1759 ();
 FILLCELL_X32 FILLCELL_144_1791 ();
 FILLCELL_X32 FILLCELL_144_1823 ();
 FILLCELL_X32 FILLCELL_144_1855 ();
 FILLCELL_X8 FILLCELL_144_1887 ();
 FILLCELL_X2 FILLCELL_144_1895 ();
 FILLCELL_X32 FILLCELL_145_0 ();
 FILLCELL_X32 FILLCELL_145_32 ();
 FILLCELL_X16 FILLCELL_145_64 ();
 FILLCELL_X2 FILLCELL_145_80 ();
 FILLCELL_X32 FILLCELL_145_85 ();
 FILLCELL_X8 FILLCELL_145_117 ();
 FILLCELL_X4 FILLCELL_145_125 ();
 FILLCELL_X2 FILLCELL_145_129 ();
 FILLCELL_X1 FILLCELL_145_131 ();
 FILLCELL_X32 FILLCELL_145_136 ();
 FILLCELL_X8 FILLCELL_145_168 ();
 FILLCELL_X2 FILLCELL_145_176 ();
 FILLCELL_X32 FILLCELL_145_181 ();
 FILLCELL_X32 FILLCELL_145_213 ();
 FILLCELL_X32 FILLCELL_145_245 ();
 FILLCELL_X8 FILLCELL_145_277 ();
 FILLCELL_X4 FILLCELL_145_285 ();
 FILLCELL_X2 FILLCELL_145_289 ();
 FILLCELL_X32 FILLCELL_145_300 ();
 FILLCELL_X32 FILLCELL_145_332 ();
 FILLCELL_X32 FILLCELL_145_364 ();
 FILLCELL_X32 FILLCELL_145_396 ();
 FILLCELL_X32 FILLCELL_145_428 ();
 FILLCELL_X8 FILLCELL_145_460 ();
 FILLCELL_X1 FILLCELL_145_468 ();
 FILLCELL_X32 FILLCELL_145_472 ();
 FILLCELL_X32 FILLCELL_145_504 ();
 FILLCELL_X32 FILLCELL_145_536 ();
 FILLCELL_X32 FILLCELL_145_568 ();
 FILLCELL_X32 FILLCELL_145_600 ();
 FILLCELL_X32 FILLCELL_145_632 ();
 FILLCELL_X32 FILLCELL_145_664 ();
 FILLCELL_X32 FILLCELL_145_696 ();
 FILLCELL_X8 FILLCELL_145_728 ();
 FILLCELL_X1 FILLCELL_145_736 ();
 FILLCELL_X32 FILLCELL_145_739 ();
 FILLCELL_X32 FILLCELL_145_771 ();
 FILLCELL_X32 FILLCELL_145_803 ();
 FILLCELL_X32 FILLCELL_145_835 ();
 FILLCELL_X32 FILLCELL_145_867 ();
 FILLCELL_X32 FILLCELL_145_899 ();
 FILLCELL_X32 FILLCELL_145_931 ();
 FILLCELL_X32 FILLCELL_145_963 ();
 FILLCELL_X32 FILLCELL_145_995 ();
 FILLCELL_X32 FILLCELL_145_1027 ();
 FILLCELL_X32 FILLCELL_145_1059 ();
 FILLCELL_X32 FILLCELL_145_1091 ();
 FILLCELL_X32 FILLCELL_145_1123 ();
 FILLCELL_X32 FILLCELL_145_1155 ();
 FILLCELL_X32 FILLCELL_145_1187 ();
 FILLCELL_X32 FILLCELL_145_1219 ();
 FILLCELL_X32 FILLCELL_145_1251 ();
 FILLCELL_X32 FILLCELL_145_1283 ();
 FILLCELL_X32 FILLCELL_145_1315 ();
 FILLCELL_X32 FILLCELL_145_1347 ();
 FILLCELL_X32 FILLCELL_145_1379 ();
 FILLCELL_X32 FILLCELL_145_1411 ();
 FILLCELL_X32 FILLCELL_145_1443 ();
 FILLCELL_X32 FILLCELL_145_1475 ();
 FILLCELL_X32 FILLCELL_145_1507 ();
 FILLCELL_X32 FILLCELL_145_1539 ();
 FILLCELL_X32 FILLCELL_145_1571 ();
 FILLCELL_X32 FILLCELL_145_1603 ();
 FILLCELL_X32 FILLCELL_145_1635 ();
 FILLCELL_X32 FILLCELL_145_1667 ();
 FILLCELL_X32 FILLCELL_145_1699 ();
 FILLCELL_X32 FILLCELL_145_1731 ();
 FILLCELL_X32 FILLCELL_145_1763 ();
 FILLCELL_X32 FILLCELL_145_1795 ();
 FILLCELL_X32 FILLCELL_145_1827 ();
 FILLCELL_X32 FILLCELL_145_1859 ();
 FILLCELL_X4 FILLCELL_145_1891 ();
 FILLCELL_X2 FILLCELL_145_1895 ();
 FILLCELL_X32 FILLCELL_146_0 ();
 FILLCELL_X32 FILLCELL_146_32 ();
 FILLCELL_X32 FILLCELL_146_64 ();
 FILLCELL_X32 FILLCELL_146_96 ();
 FILLCELL_X32 FILLCELL_146_128 ();
 FILLCELL_X32 FILLCELL_146_160 ();
 FILLCELL_X32 FILLCELL_146_192 ();
 FILLCELL_X32 FILLCELL_146_224 ();
 FILLCELL_X32 FILLCELL_146_256 ();
 FILLCELL_X32 FILLCELL_146_288 ();
 FILLCELL_X32 FILLCELL_146_320 ();
 FILLCELL_X32 FILLCELL_146_352 ();
 FILLCELL_X32 FILLCELL_146_384 ();
 FILLCELL_X32 FILLCELL_146_416 ();
 FILLCELL_X32 FILLCELL_146_448 ();
 FILLCELL_X32 FILLCELL_146_480 ();
 FILLCELL_X32 FILLCELL_146_512 ();
 FILLCELL_X16 FILLCELL_146_544 ();
 FILLCELL_X8 FILLCELL_146_560 ();
 FILLCELL_X4 FILLCELL_146_568 ();
 FILLCELL_X1 FILLCELL_146_572 ();
 FILLCELL_X32 FILLCELL_146_576 ();
 FILLCELL_X32 FILLCELL_146_608 ();
 FILLCELL_X32 FILLCELL_146_640 ();
 FILLCELL_X32 FILLCELL_146_672 ();
 FILLCELL_X16 FILLCELL_146_704 ();
 FILLCELL_X8 FILLCELL_146_720 ();
 FILLCELL_X4 FILLCELL_146_728 ();
 FILLCELL_X1 FILLCELL_146_732 ();
 FILLCELL_X32 FILLCELL_146_739 ();
 FILLCELL_X32 FILLCELL_146_771 ();
 FILLCELL_X32 FILLCELL_146_803 ();
 FILLCELL_X32 FILLCELL_146_835 ();
 FILLCELL_X32 FILLCELL_146_867 ();
 FILLCELL_X16 FILLCELL_146_899 ();
 FILLCELL_X8 FILLCELL_146_915 ();
 FILLCELL_X4 FILLCELL_146_923 ();
 FILLCELL_X2 FILLCELL_146_927 ();
 FILLCELL_X32 FILLCELL_146_933 ();
 FILLCELL_X32 FILLCELL_146_965 ();
 FILLCELL_X32 FILLCELL_146_997 ();
 FILLCELL_X32 FILLCELL_146_1029 ();
 FILLCELL_X32 FILLCELL_146_1061 ();
 FILLCELL_X32 FILLCELL_146_1093 ();
 FILLCELL_X32 FILLCELL_146_1125 ();
 FILLCELL_X32 FILLCELL_146_1157 ();
 FILLCELL_X32 FILLCELL_146_1189 ();
 FILLCELL_X32 FILLCELL_146_1221 ();
 FILLCELL_X32 FILLCELL_146_1253 ();
 FILLCELL_X32 FILLCELL_146_1285 ();
 FILLCELL_X32 FILLCELL_146_1317 ();
 FILLCELL_X32 FILLCELL_146_1349 ();
 FILLCELL_X32 FILLCELL_146_1381 ();
 FILLCELL_X32 FILLCELL_146_1413 ();
 FILLCELL_X32 FILLCELL_146_1445 ();
 FILLCELL_X32 FILLCELL_146_1477 ();
 FILLCELL_X32 FILLCELL_146_1509 ();
 FILLCELL_X32 FILLCELL_146_1541 ();
 FILLCELL_X32 FILLCELL_146_1573 ();
 FILLCELL_X32 FILLCELL_146_1605 ();
 FILLCELL_X32 FILLCELL_146_1637 ();
 FILLCELL_X32 FILLCELL_146_1669 ();
 FILLCELL_X32 FILLCELL_146_1701 ();
 FILLCELL_X32 FILLCELL_146_1733 ();
 FILLCELL_X32 FILLCELL_146_1765 ();
 FILLCELL_X32 FILLCELL_146_1797 ();
 FILLCELL_X32 FILLCELL_146_1829 ();
 FILLCELL_X32 FILLCELL_146_1861 ();
 FILLCELL_X4 FILLCELL_146_1893 ();
 FILLCELL_X32 FILLCELL_147_0 ();
 FILLCELL_X32 FILLCELL_147_32 ();
 FILLCELL_X16 FILLCELL_147_64 ();
 FILLCELL_X8 FILLCELL_147_80 ();
 FILLCELL_X4 FILLCELL_147_88 ();
 FILLCELL_X1 FILLCELL_147_92 ();
 FILLCELL_X32 FILLCELL_147_97 ();
 FILLCELL_X32 FILLCELL_147_129 ();
 FILLCELL_X32 FILLCELL_147_161 ();
 FILLCELL_X32 FILLCELL_147_193 ();
 FILLCELL_X32 FILLCELL_147_225 ();
 FILLCELL_X32 FILLCELL_147_257 ();
 FILLCELL_X32 FILLCELL_147_289 ();
 FILLCELL_X32 FILLCELL_147_321 ();
 FILLCELL_X32 FILLCELL_147_353 ();
 FILLCELL_X32 FILLCELL_147_385 ();
 FILLCELL_X32 FILLCELL_147_417 ();
 FILLCELL_X32 FILLCELL_147_449 ();
 FILLCELL_X8 FILLCELL_147_481 ();
 FILLCELL_X4 FILLCELL_147_489 ();
 FILLCELL_X1 FILLCELL_147_493 ();
 FILLCELL_X32 FILLCELL_147_498 ();
 FILLCELL_X32 FILLCELL_147_530 ();
 FILLCELL_X32 FILLCELL_147_562 ();
 FILLCELL_X32 FILLCELL_147_594 ();
 FILLCELL_X32 FILLCELL_147_626 ();
 FILLCELL_X32 FILLCELL_147_658 ();
 FILLCELL_X32 FILLCELL_147_690 ();
 FILLCELL_X32 FILLCELL_147_722 ();
 FILLCELL_X32 FILLCELL_147_754 ();
 FILLCELL_X32 FILLCELL_147_786 ();
 FILLCELL_X32 FILLCELL_147_818 ();
 FILLCELL_X32 FILLCELL_147_850 ();
 FILLCELL_X32 FILLCELL_147_882 ();
 FILLCELL_X32 FILLCELL_147_914 ();
 FILLCELL_X8 FILLCELL_147_946 ();
 FILLCELL_X32 FILLCELL_147_958 ();
 FILLCELL_X8 FILLCELL_147_990 ();
 FILLCELL_X2 FILLCELL_147_998 ();
 FILLCELL_X1 FILLCELL_147_1000 ();
 FILLCELL_X32 FILLCELL_147_1018 ();
 FILLCELL_X32 FILLCELL_147_1050 ();
 FILLCELL_X32 FILLCELL_147_1082 ();
 FILLCELL_X32 FILLCELL_147_1114 ();
 FILLCELL_X32 FILLCELL_147_1146 ();
 FILLCELL_X32 FILLCELL_147_1178 ();
 FILLCELL_X32 FILLCELL_147_1210 ();
 FILLCELL_X32 FILLCELL_147_1242 ();
 FILLCELL_X32 FILLCELL_147_1274 ();
 FILLCELL_X32 FILLCELL_147_1306 ();
 FILLCELL_X32 FILLCELL_147_1338 ();
 FILLCELL_X32 FILLCELL_147_1370 ();
 FILLCELL_X32 FILLCELL_147_1402 ();
 FILLCELL_X32 FILLCELL_147_1434 ();
 FILLCELL_X32 FILLCELL_147_1466 ();
 FILLCELL_X32 FILLCELL_147_1498 ();
 FILLCELL_X32 FILLCELL_147_1530 ();
 FILLCELL_X32 FILLCELL_147_1562 ();
 FILLCELL_X32 FILLCELL_147_1594 ();
 FILLCELL_X32 FILLCELL_147_1626 ();
 FILLCELL_X32 FILLCELL_147_1658 ();
 FILLCELL_X32 FILLCELL_147_1690 ();
 FILLCELL_X32 FILLCELL_147_1722 ();
 FILLCELL_X32 FILLCELL_147_1754 ();
 FILLCELL_X32 FILLCELL_147_1786 ();
 FILLCELL_X32 FILLCELL_147_1818 ();
 FILLCELL_X32 FILLCELL_147_1850 ();
 FILLCELL_X8 FILLCELL_147_1882 ();
 FILLCELL_X4 FILLCELL_147_1890 ();
 FILLCELL_X2 FILLCELL_147_1894 ();
 FILLCELL_X1 FILLCELL_147_1896 ();
 FILLCELL_X32 FILLCELL_148_0 ();
 FILLCELL_X32 FILLCELL_148_32 ();
 FILLCELL_X32 FILLCELL_148_64 ();
 FILLCELL_X32 FILLCELL_148_96 ();
 FILLCELL_X32 FILLCELL_148_128 ();
 FILLCELL_X32 FILLCELL_148_160 ();
 FILLCELL_X32 FILLCELL_148_192 ();
 FILLCELL_X32 FILLCELL_148_224 ();
 FILLCELL_X32 FILLCELL_148_256 ();
 FILLCELL_X32 FILLCELL_148_288 ();
 FILLCELL_X32 FILLCELL_148_320 ();
 FILLCELL_X32 FILLCELL_148_352 ();
 FILLCELL_X32 FILLCELL_148_384 ();
 FILLCELL_X32 FILLCELL_148_416 ();
 FILLCELL_X32 FILLCELL_148_448 ();
 FILLCELL_X16 FILLCELL_148_480 ();
 FILLCELL_X4 FILLCELL_148_496 ();
 FILLCELL_X1 FILLCELL_148_500 ();
 FILLCELL_X32 FILLCELL_148_503 ();
 FILLCELL_X32 FILLCELL_148_535 ();
 FILLCELL_X16 FILLCELL_148_567 ();
 FILLCELL_X8 FILLCELL_148_583 ();
 FILLCELL_X1 FILLCELL_148_591 ();
 FILLCELL_X4 FILLCELL_148_594 ();
 FILLCELL_X2 FILLCELL_148_598 ();
 FILLCELL_X32 FILLCELL_148_604 ();
 FILLCELL_X32 FILLCELL_148_636 ();
 FILLCELL_X32 FILLCELL_148_668 ();
 FILLCELL_X32 FILLCELL_148_700 ();
 FILLCELL_X32 FILLCELL_148_732 ();
 FILLCELL_X4 FILLCELL_148_764 ();
 FILLCELL_X2 FILLCELL_148_768 ();
 FILLCELL_X1 FILLCELL_148_770 ();
 FILLCELL_X32 FILLCELL_148_775 ();
 FILLCELL_X32 FILLCELL_148_807 ();
 FILLCELL_X32 FILLCELL_148_839 ();
 FILLCELL_X32 FILLCELL_148_871 ();
 FILLCELL_X32 FILLCELL_148_903 ();
 FILLCELL_X4 FILLCELL_148_935 ();
 FILLCELL_X1 FILLCELL_148_939 ();
 FILLCELL_X32 FILLCELL_148_943 ();
 FILLCELL_X32 FILLCELL_148_975 ();
 FILLCELL_X32 FILLCELL_148_1007 ();
 FILLCELL_X32 FILLCELL_148_1039 ();
 FILLCELL_X32 FILLCELL_148_1071 ();
 FILLCELL_X32 FILLCELL_148_1103 ();
 FILLCELL_X32 FILLCELL_148_1135 ();
 FILLCELL_X32 FILLCELL_148_1167 ();
 FILLCELL_X32 FILLCELL_148_1199 ();
 FILLCELL_X32 FILLCELL_148_1231 ();
 FILLCELL_X32 FILLCELL_148_1263 ();
 FILLCELL_X32 FILLCELL_148_1295 ();
 FILLCELL_X32 FILLCELL_148_1327 ();
 FILLCELL_X32 FILLCELL_148_1359 ();
 FILLCELL_X32 FILLCELL_148_1391 ();
 FILLCELL_X32 FILLCELL_148_1423 ();
 FILLCELL_X32 FILLCELL_148_1455 ();
 FILLCELL_X32 FILLCELL_148_1487 ();
 FILLCELL_X32 FILLCELL_148_1519 ();
 FILLCELL_X32 FILLCELL_148_1551 ();
 FILLCELL_X32 FILLCELL_148_1583 ();
 FILLCELL_X32 FILLCELL_148_1615 ();
 FILLCELL_X32 FILLCELL_148_1647 ();
 FILLCELL_X32 FILLCELL_148_1679 ();
 FILLCELL_X32 FILLCELL_148_1711 ();
 FILLCELL_X32 FILLCELL_148_1743 ();
 FILLCELL_X32 FILLCELL_148_1775 ();
 FILLCELL_X32 FILLCELL_148_1807 ();
 FILLCELL_X32 FILLCELL_148_1839 ();
 FILLCELL_X16 FILLCELL_148_1871 ();
 FILLCELL_X8 FILLCELL_148_1887 ();
 FILLCELL_X2 FILLCELL_148_1895 ();
 FILLCELL_X32 FILLCELL_149_0 ();
 FILLCELL_X8 FILLCELL_149_32 ();
 FILLCELL_X32 FILLCELL_149_57 ();
 FILLCELL_X32 FILLCELL_149_89 ();
 FILLCELL_X32 FILLCELL_149_121 ();
 FILLCELL_X32 FILLCELL_149_153 ();
 FILLCELL_X32 FILLCELL_149_185 ();
 FILLCELL_X32 FILLCELL_149_217 ();
 FILLCELL_X32 FILLCELL_149_249 ();
 FILLCELL_X32 FILLCELL_149_281 ();
 FILLCELL_X32 FILLCELL_149_313 ();
 FILLCELL_X32 FILLCELL_149_345 ();
 FILLCELL_X4 FILLCELL_149_377 ();
 FILLCELL_X2 FILLCELL_149_381 ();
 FILLCELL_X1 FILLCELL_149_383 ();
 FILLCELL_X32 FILLCELL_149_389 ();
 FILLCELL_X16 FILLCELL_149_421 ();
 FILLCELL_X4 FILLCELL_149_437 ();
 FILLCELL_X2 FILLCELL_149_441 ();
 FILLCELL_X32 FILLCELL_149_446 ();
 FILLCELL_X1 FILLCELL_149_478 ();
 FILLCELL_X32 FILLCELL_149_481 ();
 FILLCELL_X32 FILLCELL_149_513 ();
 FILLCELL_X32 FILLCELL_149_545 ();
 FILLCELL_X16 FILLCELL_149_577 ();
 FILLCELL_X2 FILLCELL_149_593 ();
 FILLCELL_X1 FILLCELL_149_595 ();
 FILLCELL_X16 FILLCELL_149_599 ();
 FILLCELL_X4 FILLCELL_149_615 ();
 FILLCELL_X1 FILLCELL_149_619 ();
 FILLCELL_X32 FILLCELL_149_622 ();
 FILLCELL_X2 FILLCELL_149_654 ();
 FILLCELL_X32 FILLCELL_149_660 ();
 FILLCELL_X32 FILLCELL_149_692 ();
 FILLCELL_X16 FILLCELL_149_724 ();
 FILLCELL_X8 FILLCELL_149_740 ();
 FILLCELL_X4 FILLCELL_149_748 ();
 FILLCELL_X32 FILLCELL_149_755 ();
 FILLCELL_X32 FILLCELL_149_787 ();
 FILLCELL_X32 FILLCELL_149_819 ();
 FILLCELL_X32 FILLCELL_149_851 ();
 FILLCELL_X32 FILLCELL_149_883 ();
 FILLCELL_X32 FILLCELL_149_915 ();
 FILLCELL_X32 FILLCELL_149_947 ();
 FILLCELL_X32 FILLCELL_149_979 ();
 FILLCELL_X32 FILLCELL_149_1011 ();
 FILLCELL_X32 FILLCELL_149_1043 ();
 FILLCELL_X8 FILLCELL_149_1075 ();
 FILLCELL_X2 FILLCELL_149_1083 ();
 FILLCELL_X1 FILLCELL_149_1085 ();
 FILLCELL_X32 FILLCELL_149_1090 ();
 FILLCELL_X32 FILLCELL_149_1122 ();
 FILLCELL_X32 FILLCELL_149_1154 ();
 FILLCELL_X32 FILLCELL_149_1186 ();
 FILLCELL_X32 FILLCELL_149_1218 ();
 FILLCELL_X32 FILLCELL_149_1250 ();
 FILLCELL_X32 FILLCELL_149_1282 ();
 FILLCELL_X32 FILLCELL_149_1314 ();
 FILLCELL_X32 FILLCELL_149_1346 ();
 FILLCELL_X32 FILLCELL_149_1378 ();
 FILLCELL_X32 FILLCELL_149_1410 ();
 FILLCELL_X32 FILLCELL_149_1442 ();
 FILLCELL_X32 FILLCELL_149_1474 ();
 FILLCELL_X32 FILLCELL_149_1506 ();
 FILLCELL_X32 FILLCELL_149_1538 ();
 FILLCELL_X32 FILLCELL_149_1570 ();
 FILLCELL_X32 FILLCELL_149_1602 ();
 FILLCELL_X32 FILLCELL_149_1634 ();
 FILLCELL_X32 FILLCELL_149_1666 ();
 FILLCELL_X32 FILLCELL_149_1698 ();
 FILLCELL_X32 FILLCELL_149_1730 ();
 FILLCELL_X32 FILLCELL_149_1762 ();
 FILLCELL_X32 FILLCELL_149_1794 ();
 FILLCELL_X32 FILLCELL_149_1826 ();
 FILLCELL_X32 FILLCELL_149_1858 ();
 FILLCELL_X4 FILLCELL_149_1890 ();
 FILLCELL_X2 FILLCELL_149_1894 ();
 FILLCELL_X1 FILLCELL_149_1896 ();
 FILLCELL_X32 FILLCELL_150_0 ();
 FILLCELL_X32 FILLCELL_150_32 ();
 FILLCELL_X32 FILLCELL_150_64 ();
 FILLCELL_X32 FILLCELL_150_96 ();
 FILLCELL_X16 FILLCELL_150_128 ();
 FILLCELL_X2 FILLCELL_150_144 ();
 FILLCELL_X32 FILLCELL_150_151 ();
 FILLCELL_X32 FILLCELL_150_183 ();
 FILLCELL_X32 FILLCELL_150_215 ();
 FILLCELL_X32 FILLCELL_150_247 ();
 FILLCELL_X32 FILLCELL_150_279 ();
 FILLCELL_X32 FILLCELL_150_311 ();
 FILLCELL_X32 FILLCELL_150_343 ();
 FILLCELL_X32 FILLCELL_150_375 ();
 FILLCELL_X32 FILLCELL_150_407 ();
 FILLCELL_X16 FILLCELL_150_439 ();
 FILLCELL_X8 FILLCELL_150_455 ();
 FILLCELL_X2 FILLCELL_150_463 ();
 FILLCELL_X1 FILLCELL_150_465 ();
 FILLCELL_X32 FILLCELL_150_469 ();
 FILLCELL_X32 FILLCELL_150_501 ();
 FILLCELL_X32 FILLCELL_150_533 ();
 FILLCELL_X32 FILLCELL_150_565 ();
 FILLCELL_X32 FILLCELL_150_597 ();
 FILLCELL_X32 FILLCELL_150_629 ();
 FILLCELL_X32 FILLCELL_150_661 ();
 FILLCELL_X32 FILLCELL_150_697 ();
 FILLCELL_X32 FILLCELL_150_729 ();
 FILLCELL_X32 FILLCELL_150_761 ();
 FILLCELL_X32 FILLCELL_150_793 ();
 FILLCELL_X32 FILLCELL_150_825 ();
 FILLCELL_X32 FILLCELL_150_857 ();
 FILLCELL_X32 FILLCELL_150_889 ();
 FILLCELL_X32 FILLCELL_150_921 ();
 FILLCELL_X32 FILLCELL_150_953 ();
 FILLCELL_X32 FILLCELL_150_985 ();
 FILLCELL_X32 FILLCELL_150_1017 ();
 FILLCELL_X32 FILLCELL_150_1049 ();
 FILLCELL_X32 FILLCELL_150_1081 ();
 FILLCELL_X32 FILLCELL_150_1113 ();
 FILLCELL_X32 FILLCELL_150_1145 ();
 FILLCELL_X32 FILLCELL_150_1177 ();
 FILLCELL_X32 FILLCELL_150_1209 ();
 FILLCELL_X32 FILLCELL_150_1241 ();
 FILLCELL_X32 FILLCELL_150_1273 ();
 FILLCELL_X32 FILLCELL_150_1305 ();
 FILLCELL_X32 FILLCELL_150_1337 ();
 FILLCELL_X32 FILLCELL_150_1369 ();
 FILLCELL_X32 FILLCELL_150_1401 ();
 FILLCELL_X32 FILLCELL_150_1433 ();
 FILLCELL_X32 FILLCELL_150_1465 ();
 FILLCELL_X32 FILLCELL_150_1497 ();
 FILLCELL_X32 FILLCELL_150_1529 ();
 FILLCELL_X32 FILLCELL_150_1561 ();
 FILLCELL_X32 FILLCELL_150_1593 ();
 FILLCELL_X32 FILLCELL_150_1625 ();
 FILLCELL_X32 FILLCELL_150_1657 ();
 FILLCELL_X32 FILLCELL_150_1689 ();
 FILLCELL_X32 FILLCELL_150_1721 ();
 FILLCELL_X32 FILLCELL_150_1753 ();
 FILLCELL_X32 FILLCELL_150_1785 ();
 FILLCELL_X32 FILLCELL_150_1817 ();
 FILLCELL_X32 FILLCELL_150_1849 ();
 FILLCELL_X16 FILLCELL_150_1881 ();
 FILLCELL_X32 FILLCELL_151_0 ();
 FILLCELL_X32 FILLCELL_151_32 ();
 FILLCELL_X32 FILLCELL_151_64 ();
 FILLCELL_X32 FILLCELL_151_96 ();
 FILLCELL_X32 FILLCELL_151_128 ();
 FILLCELL_X4 FILLCELL_151_160 ();
 FILLCELL_X1 FILLCELL_151_164 ();
 FILLCELL_X32 FILLCELL_151_167 ();
 FILLCELL_X16 FILLCELL_151_199 ();
 FILLCELL_X8 FILLCELL_151_215 ();
 FILLCELL_X4 FILLCELL_151_223 ();
 FILLCELL_X1 FILLCELL_151_227 ();
 FILLCELL_X16 FILLCELL_151_246 ();
 FILLCELL_X8 FILLCELL_151_262 ();
 FILLCELL_X4 FILLCELL_151_270 ();
 FILLCELL_X2 FILLCELL_151_274 ();
 FILLCELL_X32 FILLCELL_151_284 ();
 FILLCELL_X32 FILLCELL_151_316 ();
 FILLCELL_X32 FILLCELL_151_348 ();
 FILLCELL_X32 FILLCELL_151_380 ();
 FILLCELL_X32 FILLCELL_151_412 ();
 FILLCELL_X32 FILLCELL_151_444 ();
 FILLCELL_X32 FILLCELL_151_476 ();
 FILLCELL_X32 FILLCELL_151_508 ();
 FILLCELL_X32 FILLCELL_151_540 ();
 FILLCELL_X32 FILLCELL_151_572 ();
 FILLCELL_X32 FILLCELL_151_604 ();
 FILLCELL_X32 FILLCELL_151_636 ();
 FILLCELL_X32 FILLCELL_151_668 ();
 FILLCELL_X16 FILLCELL_151_700 ();
 FILLCELL_X8 FILLCELL_151_716 ();
 FILLCELL_X4 FILLCELL_151_724 ();
 FILLCELL_X2 FILLCELL_151_728 ();
 FILLCELL_X1 FILLCELL_151_730 ();
 FILLCELL_X32 FILLCELL_151_734 ();
 FILLCELL_X16 FILLCELL_151_766 ();
 FILLCELL_X8 FILLCELL_151_782 ();
 FILLCELL_X2 FILLCELL_151_790 ();
 FILLCELL_X4 FILLCELL_151_797 ();
 FILLCELL_X32 FILLCELL_151_803 ();
 FILLCELL_X32 FILLCELL_151_835 ();
 FILLCELL_X32 FILLCELL_151_867 ();
 FILLCELL_X32 FILLCELL_151_899 ();
 FILLCELL_X32 FILLCELL_151_931 ();
 FILLCELL_X32 FILLCELL_151_963 ();
 FILLCELL_X32 FILLCELL_151_995 ();
 FILLCELL_X32 FILLCELL_151_1027 ();
 FILLCELL_X32 FILLCELL_151_1059 ();
 FILLCELL_X2 FILLCELL_151_1091 ();
 FILLCELL_X32 FILLCELL_151_1098 ();
 FILLCELL_X32 FILLCELL_151_1130 ();
 FILLCELL_X32 FILLCELL_151_1162 ();
 FILLCELL_X32 FILLCELL_151_1194 ();
 FILLCELL_X32 FILLCELL_151_1226 ();
 FILLCELL_X32 FILLCELL_151_1258 ();
 FILLCELL_X32 FILLCELL_151_1290 ();
 FILLCELL_X32 FILLCELL_151_1322 ();
 FILLCELL_X32 FILLCELL_151_1354 ();
 FILLCELL_X32 FILLCELL_151_1386 ();
 FILLCELL_X32 FILLCELL_151_1418 ();
 FILLCELL_X32 FILLCELL_151_1450 ();
 FILLCELL_X32 FILLCELL_151_1482 ();
 FILLCELL_X32 FILLCELL_151_1514 ();
 FILLCELL_X32 FILLCELL_151_1546 ();
 FILLCELL_X32 FILLCELL_151_1578 ();
 FILLCELL_X32 FILLCELL_151_1610 ();
 FILLCELL_X32 FILLCELL_151_1642 ();
 FILLCELL_X32 FILLCELL_151_1674 ();
 FILLCELL_X32 FILLCELL_151_1706 ();
 FILLCELL_X32 FILLCELL_151_1738 ();
 FILLCELL_X32 FILLCELL_151_1770 ();
 FILLCELL_X32 FILLCELL_151_1802 ();
 FILLCELL_X32 FILLCELL_151_1834 ();
 FILLCELL_X16 FILLCELL_151_1866 ();
 FILLCELL_X8 FILLCELL_151_1882 ();
 FILLCELL_X4 FILLCELL_151_1890 ();
 FILLCELL_X2 FILLCELL_151_1894 ();
 FILLCELL_X1 FILLCELL_151_1896 ();
 FILLCELL_X32 FILLCELL_152_0 ();
 FILLCELL_X32 FILLCELL_152_32 ();
 FILLCELL_X32 FILLCELL_152_64 ();
 FILLCELL_X32 FILLCELL_152_96 ();
 FILLCELL_X32 FILLCELL_152_128 ();
 FILLCELL_X32 FILLCELL_152_164 ();
 FILLCELL_X32 FILLCELL_152_196 ();
 FILLCELL_X32 FILLCELL_152_228 ();
 FILLCELL_X32 FILLCELL_152_260 ();
 FILLCELL_X32 FILLCELL_152_292 ();
 FILLCELL_X32 FILLCELL_152_324 ();
 FILLCELL_X8 FILLCELL_152_356 ();
 FILLCELL_X4 FILLCELL_152_364 ();
 FILLCELL_X2 FILLCELL_152_368 ();
 FILLCELL_X1 FILLCELL_152_370 ();
 FILLCELL_X32 FILLCELL_152_380 ();
 FILLCELL_X32 FILLCELL_152_412 ();
 FILLCELL_X32 FILLCELL_152_444 ();
 FILLCELL_X32 FILLCELL_152_476 ();
 FILLCELL_X32 FILLCELL_152_508 ();
 FILLCELL_X32 FILLCELL_152_540 ();
 FILLCELL_X16 FILLCELL_152_572 ();
 FILLCELL_X4 FILLCELL_152_588 ();
 FILLCELL_X2 FILLCELL_152_592 ();
 FILLCELL_X32 FILLCELL_152_598 ();
 FILLCELL_X32 FILLCELL_152_630 ();
 FILLCELL_X32 FILLCELL_152_662 ();
 FILLCELL_X32 FILLCELL_152_694 ();
 FILLCELL_X32 FILLCELL_152_726 ();
 FILLCELL_X32 FILLCELL_152_758 ();
 FILLCELL_X32 FILLCELL_152_790 ();
 FILLCELL_X32 FILLCELL_152_822 ();
 FILLCELL_X32 FILLCELL_152_854 ();
 FILLCELL_X32 FILLCELL_152_886 ();
 FILLCELL_X32 FILLCELL_152_918 ();
 FILLCELL_X32 FILLCELL_152_950 ();
 FILLCELL_X32 FILLCELL_152_982 ();
 FILLCELL_X32 FILLCELL_152_1014 ();
 FILLCELL_X32 FILLCELL_152_1046 ();
 FILLCELL_X32 FILLCELL_152_1078 ();
 FILLCELL_X32 FILLCELL_152_1110 ();
 FILLCELL_X32 FILLCELL_152_1142 ();
 FILLCELL_X32 FILLCELL_152_1174 ();
 FILLCELL_X32 FILLCELL_152_1206 ();
 FILLCELL_X32 FILLCELL_152_1238 ();
 FILLCELL_X32 FILLCELL_152_1270 ();
 FILLCELL_X32 FILLCELL_152_1302 ();
 FILLCELL_X32 FILLCELL_152_1334 ();
 FILLCELL_X32 FILLCELL_152_1366 ();
 FILLCELL_X32 FILLCELL_152_1398 ();
 FILLCELL_X32 FILLCELL_152_1430 ();
 FILLCELL_X32 FILLCELL_152_1462 ();
 FILLCELL_X32 FILLCELL_152_1494 ();
 FILLCELL_X32 FILLCELL_152_1526 ();
 FILLCELL_X32 FILLCELL_152_1558 ();
 FILLCELL_X32 FILLCELL_152_1590 ();
 FILLCELL_X32 FILLCELL_152_1622 ();
 FILLCELL_X32 FILLCELL_152_1654 ();
 FILLCELL_X32 FILLCELL_152_1686 ();
 FILLCELL_X32 FILLCELL_152_1718 ();
 FILLCELL_X32 FILLCELL_152_1750 ();
 FILLCELL_X32 FILLCELL_152_1782 ();
 FILLCELL_X32 FILLCELL_152_1814 ();
 FILLCELL_X32 FILLCELL_152_1846 ();
 FILLCELL_X16 FILLCELL_152_1878 ();
 FILLCELL_X2 FILLCELL_152_1894 ();
 FILLCELL_X1 FILLCELL_152_1896 ();
 FILLCELL_X32 FILLCELL_153_0 ();
 FILLCELL_X32 FILLCELL_153_32 ();
 FILLCELL_X32 FILLCELL_153_64 ();
 FILLCELL_X32 FILLCELL_153_96 ();
 FILLCELL_X32 FILLCELL_153_128 ();
 FILLCELL_X32 FILLCELL_153_160 ();
 FILLCELL_X32 FILLCELL_153_192 ();
 FILLCELL_X32 FILLCELL_153_224 ();
 FILLCELL_X32 FILLCELL_153_256 ();
 FILLCELL_X32 FILLCELL_153_288 ();
 FILLCELL_X32 FILLCELL_153_320 ();
 FILLCELL_X32 FILLCELL_153_352 ();
 FILLCELL_X32 FILLCELL_153_384 ();
 FILLCELL_X32 FILLCELL_153_416 ();
 FILLCELL_X32 FILLCELL_153_448 ();
 FILLCELL_X8 FILLCELL_153_480 ();
 FILLCELL_X4 FILLCELL_153_488 ();
 FILLCELL_X1 FILLCELL_153_492 ();
 FILLCELL_X32 FILLCELL_153_498 ();
 FILLCELL_X32 FILLCELL_153_530 ();
 FILLCELL_X32 FILLCELL_153_562 ();
 FILLCELL_X32 FILLCELL_153_594 ();
 FILLCELL_X32 FILLCELL_153_626 ();
 FILLCELL_X16 FILLCELL_153_658 ();
 FILLCELL_X32 FILLCELL_153_677 ();
 FILLCELL_X32 FILLCELL_153_709 ();
 FILLCELL_X32 FILLCELL_153_741 ();
 FILLCELL_X32 FILLCELL_153_773 ();
 FILLCELL_X32 FILLCELL_153_805 ();
 FILLCELL_X16 FILLCELL_153_837 ();
 FILLCELL_X2 FILLCELL_153_853 ();
 FILLCELL_X32 FILLCELL_153_861 ();
 FILLCELL_X32 FILLCELL_153_893 ();
 FILLCELL_X32 FILLCELL_153_925 ();
 FILLCELL_X32 FILLCELL_153_957 ();
 FILLCELL_X32 FILLCELL_153_989 ();
 FILLCELL_X32 FILLCELL_153_1021 ();
 FILLCELL_X32 FILLCELL_153_1053 ();
 FILLCELL_X32 FILLCELL_153_1085 ();
 FILLCELL_X32 FILLCELL_153_1117 ();
 FILLCELL_X32 FILLCELL_153_1149 ();
 FILLCELL_X32 FILLCELL_153_1181 ();
 FILLCELL_X32 FILLCELL_153_1213 ();
 FILLCELL_X32 FILLCELL_153_1245 ();
 FILLCELL_X32 FILLCELL_153_1277 ();
 FILLCELL_X32 FILLCELL_153_1309 ();
 FILLCELL_X32 FILLCELL_153_1341 ();
 FILLCELL_X32 FILLCELL_153_1373 ();
 FILLCELL_X32 FILLCELL_153_1405 ();
 FILLCELL_X32 FILLCELL_153_1437 ();
 FILLCELL_X32 FILLCELL_153_1469 ();
 FILLCELL_X32 FILLCELL_153_1501 ();
 FILLCELL_X32 FILLCELL_153_1533 ();
 FILLCELL_X32 FILLCELL_153_1565 ();
 FILLCELL_X32 FILLCELL_153_1597 ();
 FILLCELL_X32 FILLCELL_153_1629 ();
 FILLCELL_X32 FILLCELL_153_1661 ();
 FILLCELL_X32 FILLCELL_153_1693 ();
 FILLCELL_X32 FILLCELL_153_1725 ();
 FILLCELL_X32 FILLCELL_153_1757 ();
 FILLCELL_X32 FILLCELL_153_1789 ();
 FILLCELL_X32 FILLCELL_153_1821 ();
 FILLCELL_X32 FILLCELL_153_1853 ();
 FILLCELL_X8 FILLCELL_153_1885 ();
 FILLCELL_X4 FILLCELL_153_1893 ();
 FILLCELL_X32 FILLCELL_154_0 ();
 FILLCELL_X32 FILLCELL_154_32 ();
 FILLCELL_X32 FILLCELL_154_64 ();
 FILLCELL_X32 FILLCELL_154_96 ();
 FILLCELL_X32 FILLCELL_154_128 ();
 FILLCELL_X32 FILLCELL_154_160 ();
 FILLCELL_X32 FILLCELL_154_192 ();
 FILLCELL_X32 FILLCELL_154_224 ();
 FILLCELL_X16 FILLCELL_154_256 ();
 FILLCELL_X8 FILLCELL_154_272 ();
 FILLCELL_X1 FILLCELL_154_280 ();
 FILLCELL_X32 FILLCELL_154_284 ();
 FILLCELL_X32 FILLCELL_154_316 ();
 FILLCELL_X32 FILLCELL_154_348 ();
 FILLCELL_X32 FILLCELL_154_380 ();
 FILLCELL_X32 FILLCELL_154_412 ();
 FILLCELL_X8 FILLCELL_154_444 ();
 FILLCELL_X32 FILLCELL_154_457 ();
 FILLCELL_X32 FILLCELL_154_489 ();
 FILLCELL_X32 FILLCELL_154_521 ();
 FILLCELL_X32 FILLCELL_154_553 ();
 FILLCELL_X32 FILLCELL_154_585 ();
 FILLCELL_X32 FILLCELL_154_617 ();
 FILLCELL_X32 FILLCELL_154_649 ();
 FILLCELL_X32 FILLCELL_154_681 ();
 FILLCELL_X32 FILLCELL_154_713 ();
 FILLCELL_X32 FILLCELL_154_745 ();
 FILLCELL_X32 FILLCELL_154_777 ();
 FILLCELL_X32 FILLCELL_154_809 ();
 FILLCELL_X32 FILLCELL_154_841 ();
 FILLCELL_X32 FILLCELL_154_873 ();
 FILLCELL_X32 FILLCELL_154_905 ();
 FILLCELL_X32 FILLCELL_154_937 ();
 FILLCELL_X32 FILLCELL_154_969 ();
 FILLCELL_X32 FILLCELL_154_1001 ();
 FILLCELL_X8 FILLCELL_154_1033 ();
 FILLCELL_X4 FILLCELL_154_1041 ();
 FILLCELL_X32 FILLCELL_154_1047 ();
 FILLCELL_X32 FILLCELL_154_1079 ();
 FILLCELL_X32 FILLCELL_154_1111 ();
 FILLCELL_X32 FILLCELL_154_1143 ();
 FILLCELL_X32 FILLCELL_154_1175 ();
 FILLCELL_X32 FILLCELL_154_1207 ();
 FILLCELL_X32 FILLCELL_154_1239 ();
 FILLCELL_X32 FILLCELL_154_1271 ();
 FILLCELL_X32 FILLCELL_154_1303 ();
 FILLCELL_X32 FILLCELL_154_1335 ();
 FILLCELL_X32 FILLCELL_154_1367 ();
 FILLCELL_X32 FILLCELL_154_1399 ();
 FILLCELL_X32 FILLCELL_154_1431 ();
 FILLCELL_X32 FILLCELL_154_1463 ();
 FILLCELL_X32 FILLCELL_154_1495 ();
 FILLCELL_X32 FILLCELL_154_1527 ();
 FILLCELL_X32 FILLCELL_154_1559 ();
 FILLCELL_X32 FILLCELL_154_1591 ();
 FILLCELL_X32 FILLCELL_154_1623 ();
 FILLCELL_X32 FILLCELL_154_1655 ();
 FILLCELL_X32 FILLCELL_154_1687 ();
 FILLCELL_X32 FILLCELL_154_1719 ();
 FILLCELL_X32 FILLCELL_154_1751 ();
 FILLCELL_X32 FILLCELL_154_1783 ();
 FILLCELL_X32 FILLCELL_154_1815 ();
 FILLCELL_X32 FILLCELL_154_1847 ();
 FILLCELL_X16 FILLCELL_154_1879 ();
 FILLCELL_X2 FILLCELL_154_1895 ();
 FILLCELL_X32 FILLCELL_155_0 ();
 FILLCELL_X32 FILLCELL_155_32 ();
 FILLCELL_X32 FILLCELL_155_64 ();
 FILLCELL_X32 FILLCELL_155_96 ();
 FILLCELL_X32 FILLCELL_155_128 ();
 FILLCELL_X16 FILLCELL_155_160 ();
 FILLCELL_X2 FILLCELL_155_176 ();
 FILLCELL_X1 FILLCELL_155_178 ();
 FILLCELL_X32 FILLCELL_155_182 ();
 FILLCELL_X32 FILLCELL_155_214 ();
 FILLCELL_X32 FILLCELL_155_246 ();
 FILLCELL_X32 FILLCELL_155_278 ();
 FILLCELL_X32 FILLCELL_155_310 ();
 FILLCELL_X32 FILLCELL_155_342 ();
 FILLCELL_X32 FILLCELL_155_374 ();
 FILLCELL_X32 FILLCELL_155_406 ();
 FILLCELL_X32 FILLCELL_155_438 ();
 FILLCELL_X32 FILLCELL_155_470 ();
 FILLCELL_X32 FILLCELL_155_502 ();
 FILLCELL_X32 FILLCELL_155_534 ();
 FILLCELL_X32 FILLCELL_155_566 ();
 FILLCELL_X32 FILLCELL_155_598 ();
 FILLCELL_X4 FILLCELL_155_630 ();
 FILLCELL_X1 FILLCELL_155_634 ();
 FILLCELL_X32 FILLCELL_155_640 ();
 FILLCELL_X32 FILLCELL_155_672 ();
 FILLCELL_X32 FILLCELL_155_704 ();
 FILLCELL_X32 FILLCELL_155_736 ();
 FILLCELL_X32 FILLCELL_155_768 ();
 FILLCELL_X32 FILLCELL_155_800 ();
 FILLCELL_X32 FILLCELL_155_832 ();
 FILLCELL_X8 FILLCELL_155_864 ();
 FILLCELL_X4 FILLCELL_155_872 ();
 FILLCELL_X16 FILLCELL_155_881 ();
 FILLCELL_X8 FILLCELL_155_897 ();
 FILLCELL_X32 FILLCELL_155_911 ();
 FILLCELL_X32 FILLCELL_155_943 ();
 FILLCELL_X32 FILLCELL_155_975 ();
 FILLCELL_X32 FILLCELL_155_1007 ();
 FILLCELL_X32 FILLCELL_155_1039 ();
 FILLCELL_X32 FILLCELL_155_1071 ();
 FILLCELL_X8 FILLCELL_155_1103 ();
 FILLCELL_X4 FILLCELL_155_1111 ();
 FILLCELL_X32 FILLCELL_155_1122 ();
 FILLCELL_X32 FILLCELL_155_1154 ();
 FILLCELL_X32 FILLCELL_155_1186 ();
 FILLCELL_X32 FILLCELL_155_1218 ();
 FILLCELL_X32 FILLCELL_155_1250 ();
 FILLCELL_X32 FILLCELL_155_1282 ();
 FILLCELL_X32 FILLCELL_155_1314 ();
 FILLCELL_X32 FILLCELL_155_1346 ();
 FILLCELL_X32 FILLCELL_155_1378 ();
 FILLCELL_X32 FILLCELL_155_1410 ();
 FILLCELL_X32 FILLCELL_155_1442 ();
 FILLCELL_X32 FILLCELL_155_1474 ();
 FILLCELL_X32 FILLCELL_155_1506 ();
 FILLCELL_X32 FILLCELL_155_1538 ();
 FILLCELL_X32 FILLCELL_155_1570 ();
 FILLCELL_X32 FILLCELL_155_1602 ();
 FILLCELL_X32 FILLCELL_155_1634 ();
 FILLCELL_X32 FILLCELL_155_1666 ();
 FILLCELL_X32 FILLCELL_155_1698 ();
 FILLCELL_X32 FILLCELL_155_1730 ();
 FILLCELL_X32 FILLCELL_155_1762 ();
 FILLCELL_X32 FILLCELL_155_1794 ();
 FILLCELL_X32 FILLCELL_155_1826 ();
 FILLCELL_X32 FILLCELL_155_1858 ();
 FILLCELL_X4 FILLCELL_155_1890 ();
 FILLCELL_X2 FILLCELL_155_1894 ();
 FILLCELL_X1 FILLCELL_155_1896 ();
 FILLCELL_X32 FILLCELL_156_0 ();
 FILLCELL_X32 FILLCELL_156_32 ();
 FILLCELL_X32 FILLCELL_156_64 ();
 FILLCELL_X32 FILLCELL_156_96 ();
 FILLCELL_X32 FILLCELL_156_128 ();
 FILLCELL_X32 FILLCELL_156_160 ();
 FILLCELL_X32 FILLCELL_156_192 ();
 FILLCELL_X32 FILLCELL_156_224 ();
 FILLCELL_X32 FILLCELL_156_256 ();
 FILLCELL_X32 FILLCELL_156_288 ();
 FILLCELL_X32 FILLCELL_156_320 ();
 FILLCELL_X32 FILLCELL_156_352 ();
 FILLCELL_X32 FILLCELL_156_384 ();
 FILLCELL_X32 FILLCELL_156_416 ();
 FILLCELL_X32 FILLCELL_156_448 ();
 FILLCELL_X32 FILLCELL_156_480 ();
 FILLCELL_X32 FILLCELL_156_512 ();
 FILLCELL_X32 FILLCELL_156_544 ();
 FILLCELL_X32 FILLCELL_156_576 ();
 FILLCELL_X32 FILLCELL_156_608 ();
 FILLCELL_X32 FILLCELL_156_640 ();
 FILLCELL_X32 FILLCELL_156_672 ();
 FILLCELL_X32 FILLCELL_156_704 ();
 FILLCELL_X32 FILLCELL_156_736 ();
 FILLCELL_X16 FILLCELL_156_768 ();
 FILLCELL_X4 FILLCELL_156_784 ();
 FILLCELL_X2 FILLCELL_156_788 ();
 FILLCELL_X32 FILLCELL_156_793 ();
 FILLCELL_X32 FILLCELL_156_825 ();
 FILLCELL_X32 FILLCELL_156_857 ();
 FILLCELL_X32 FILLCELL_156_889 ();
 FILLCELL_X32 FILLCELL_156_921 ();
 FILLCELL_X32 FILLCELL_156_953 ();
 FILLCELL_X32 FILLCELL_156_985 ();
 FILLCELL_X32 FILLCELL_156_1017 ();
 FILLCELL_X32 FILLCELL_156_1049 ();
 FILLCELL_X32 FILLCELL_156_1081 ();
 FILLCELL_X32 FILLCELL_156_1113 ();
 FILLCELL_X32 FILLCELL_156_1145 ();
 FILLCELL_X32 FILLCELL_156_1194 ();
 FILLCELL_X32 FILLCELL_156_1226 ();
 FILLCELL_X32 FILLCELL_156_1258 ();
 FILLCELL_X32 FILLCELL_156_1290 ();
 FILLCELL_X32 FILLCELL_156_1322 ();
 FILLCELL_X32 FILLCELL_156_1354 ();
 FILLCELL_X32 FILLCELL_156_1386 ();
 FILLCELL_X32 FILLCELL_156_1418 ();
 FILLCELL_X32 FILLCELL_156_1450 ();
 FILLCELL_X32 FILLCELL_156_1482 ();
 FILLCELL_X32 FILLCELL_156_1514 ();
 FILLCELL_X32 FILLCELL_156_1546 ();
 FILLCELL_X32 FILLCELL_156_1578 ();
 FILLCELL_X32 FILLCELL_156_1610 ();
 FILLCELL_X32 FILLCELL_156_1642 ();
 FILLCELL_X32 FILLCELL_156_1674 ();
 FILLCELL_X32 FILLCELL_156_1706 ();
 FILLCELL_X32 FILLCELL_156_1738 ();
 FILLCELL_X32 FILLCELL_156_1770 ();
 FILLCELL_X32 FILLCELL_156_1802 ();
 FILLCELL_X32 FILLCELL_156_1834 ();
 FILLCELL_X16 FILLCELL_156_1866 ();
 FILLCELL_X8 FILLCELL_156_1882 ();
 FILLCELL_X4 FILLCELL_156_1890 ();
 FILLCELL_X2 FILLCELL_156_1894 ();
 FILLCELL_X1 FILLCELL_156_1896 ();
 FILLCELL_X32 FILLCELL_157_0 ();
 FILLCELL_X32 FILLCELL_157_32 ();
 FILLCELL_X32 FILLCELL_157_64 ();
 FILLCELL_X32 FILLCELL_157_96 ();
 FILLCELL_X32 FILLCELL_157_128 ();
 FILLCELL_X32 FILLCELL_157_160 ();
 FILLCELL_X32 FILLCELL_157_192 ();
 FILLCELL_X32 FILLCELL_157_224 ();
 FILLCELL_X32 FILLCELL_157_256 ();
 FILLCELL_X32 FILLCELL_157_288 ();
 FILLCELL_X8 FILLCELL_157_320 ();
 FILLCELL_X32 FILLCELL_157_334 ();
 FILLCELL_X32 FILLCELL_157_366 ();
 FILLCELL_X32 FILLCELL_157_398 ();
 FILLCELL_X32 FILLCELL_157_430 ();
 FILLCELL_X32 FILLCELL_157_462 ();
 FILLCELL_X32 FILLCELL_157_494 ();
 FILLCELL_X16 FILLCELL_157_526 ();
 FILLCELL_X8 FILLCELL_157_542 ();
 FILLCELL_X32 FILLCELL_157_555 ();
 FILLCELL_X32 FILLCELL_157_587 ();
 FILLCELL_X32 FILLCELL_157_619 ();
 FILLCELL_X32 FILLCELL_157_651 ();
 FILLCELL_X32 FILLCELL_157_683 ();
 FILLCELL_X32 FILLCELL_157_715 ();
 FILLCELL_X16 FILLCELL_157_747 ();
 FILLCELL_X2 FILLCELL_157_763 ();
 FILLCELL_X1 FILLCELL_157_765 ();
 FILLCELL_X32 FILLCELL_157_768 ();
 FILLCELL_X32 FILLCELL_157_800 ();
 FILLCELL_X32 FILLCELL_157_832 ();
 FILLCELL_X32 FILLCELL_157_864 ();
 FILLCELL_X32 FILLCELL_157_896 ();
 FILLCELL_X32 FILLCELL_157_928 ();
 FILLCELL_X32 FILLCELL_157_960 ();
 FILLCELL_X32 FILLCELL_157_992 ();
 FILLCELL_X32 FILLCELL_157_1024 ();
 FILLCELL_X32 FILLCELL_157_1056 ();
 FILLCELL_X32 FILLCELL_157_1088 ();
 FILLCELL_X32 FILLCELL_157_1120 ();
 FILLCELL_X32 FILLCELL_157_1152 ();
 FILLCELL_X32 FILLCELL_157_1184 ();
 FILLCELL_X32 FILLCELL_157_1216 ();
 FILLCELL_X32 FILLCELL_157_1248 ();
 FILLCELL_X32 FILLCELL_157_1280 ();
 FILLCELL_X32 FILLCELL_157_1312 ();
 FILLCELL_X32 FILLCELL_157_1344 ();
 FILLCELL_X32 FILLCELL_157_1376 ();
 FILLCELL_X32 FILLCELL_157_1408 ();
 FILLCELL_X32 FILLCELL_157_1440 ();
 FILLCELL_X32 FILLCELL_157_1472 ();
 FILLCELL_X32 FILLCELL_157_1504 ();
 FILLCELL_X32 FILLCELL_157_1536 ();
 FILLCELL_X32 FILLCELL_157_1568 ();
 FILLCELL_X32 FILLCELL_157_1600 ();
 FILLCELL_X32 FILLCELL_157_1632 ();
 FILLCELL_X32 FILLCELL_157_1664 ();
 FILLCELL_X32 FILLCELL_157_1696 ();
 FILLCELL_X32 FILLCELL_157_1728 ();
 FILLCELL_X32 FILLCELL_157_1760 ();
 FILLCELL_X32 FILLCELL_157_1792 ();
 FILLCELL_X32 FILLCELL_157_1824 ();
 FILLCELL_X32 FILLCELL_157_1856 ();
 FILLCELL_X8 FILLCELL_157_1888 ();
 FILLCELL_X1 FILLCELL_157_1896 ();
 FILLCELL_X32 FILLCELL_158_0 ();
 FILLCELL_X32 FILLCELL_158_32 ();
 FILLCELL_X32 FILLCELL_158_64 ();
 FILLCELL_X32 FILLCELL_158_96 ();
 FILLCELL_X32 FILLCELL_158_128 ();
 FILLCELL_X32 FILLCELL_158_160 ();
 FILLCELL_X32 FILLCELL_158_192 ();
 FILLCELL_X32 FILLCELL_158_224 ();
 FILLCELL_X32 FILLCELL_158_256 ();
 FILLCELL_X8 FILLCELL_158_288 ();
 FILLCELL_X2 FILLCELL_158_296 ();
 FILLCELL_X1 FILLCELL_158_298 ();
 FILLCELL_X32 FILLCELL_158_302 ();
 FILLCELL_X32 FILLCELL_158_334 ();
 FILLCELL_X32 FILLCELL_158_366 ();
 FILLCELL_X32 FILLCELL_158_398 ();
 FILLCELL_X32 FILLCELL_158_430 ();
 FILLCELL_X32 FILLCELL_158_462 ();
 FILLCELL_X32 FILLCELL_158_494 ();
 FILLCELL_X32 FILLCELL_158_526 ();
 FILLCELL_X32 FILLCELL_158_558 ();
 FILLCELL_X32 FILLCELL_158_590 ();
 FILLCELL_X32 FILLCELL_158_622 ();
 FILLCELL_X32 FILLCELL_158_654 ();
 FILLCELL_X32 FILLCELL_158_686 ();
 FILLCELL_X32 FILLCELL_158_718 ();
 FILLCELL_X8 FILLCELL_158_750 ();
 FILLCELL_X4 FILLCELL_158_758 ();
 FILLCELL_X32 FILLCELL_158_765 ();
 FILLCELL_X32 FILLCELL_158_797 ();
 FILLCELL_X32 FILLCELL_158_829 ();
 FILLCELL_X16 FILLCELL_158_861 ();
 FILLCELL_X8 FILLCELL_158_877 ();
 FILLCELL_X4 FILLCELL_158_885 ();
 FILLCELL_X1 FILLCELL_158_889 ();
 FILLCELL_X32 FILLCELL_158_895 ();
 FILLCELL_X32 FILLCELL_158_927 ();
 FILLCELL_X32 FILLCELL_158_959 ();
 FILLCELL_X1 FILLCELL_158_991 ();
 FILLCELL_X32 FILLCELL_158_997 ();
 FILLCELL_X32 FILLCELL_158_1029 ();
 FILLCELL_X8 FILLCELL_158_1061 ();
 FILLCELL_X16 FILLCELL_158_1074 ();
 FILLCELL_X8 FILLCELL_158_1090 ();
 FILLCELL_X4 FILLCELL_158_1098 ();
 FILLCELL_X1 FILLCELL_158_1102 ();
 FILLCELL_X32 FILLCELL_158_1106 ();
 FILLCELL_X32 FILLCELL_158_1138 ();
 FILLCELL_X32 FILLCELL_158_1170 ();
 FILLCELL_X32 FILLCELL_158_1202 ();
 FILLCELL_X32 FILLCELL_158_1234 ();
 FILLCELL_X32 FILLCELL_158_1266 ();
 FILLCELL_X32 FILLCELL_158_1298 ();
 FILLCELL_X32 FILLCELL_158_1330 ();
 FILLCELL_X32 FILLCELL_158_1362 ();
 FILLCELL_X32 FILLCELL_158_1394 ();
 FILLCELL_X32 FILLCELL_158_1426 ();
 FILLCELL_X32 FILLCELL_158_1458 ();
 FILLCELL_X32 FILLCELL_158_1490 ();
 FILLCELL_X32 FILLCELL_158_1522 ();
 FILLCELL_X32 FILLCELL_158_1554 ();
 FILLCELL_X32 FILLCELL_158_1586 ();
 FILLCELL_X32 FILLCELL_158_1618 ();
 FILLCELL_X32 FILLCELL_158_1650 ();
 FILLCELL_X32 FILLCELL_158_1682 ();
 FILLCELL_X32 FILLCELL_158_1714 ();
 FILLCELL_X32 FILLCELL_158_1746 ();
 FILLCELL_X32 FILLCELL_158_1778 ();
 FILLCELL_X32 FILLCELL_158_1810 ();
 FILLCELL_X32 FILLCELL_158_1842 ();
 FILLCELL_X16 FILLCELL_158_1874 ();
 FILLCELL_X4 FILLCELL_158_1890 ();
 FILLCELL_X2 FILLCELL_158_1894 ();
 FILLCELL_X1 FILLCELL_158_1896 ();
 FILLCELL_X32 FILLCELL_159_0 ();
 FILLCELL_X32 FILLCELL_159_32 ();
 FILLCELL_X32 FILLCELL_159_64 ();
 FILLCELL_X32 FILLCELL_159_96 ();
 FILLCELL_X32 FILLCELL_159_128 ();
 FILLCELL_X32 FILLCELL_159_160 ();
 FILLCELL_X32 FILLCELL_159_192 ();
 FILLCELL_X32 FILLCELL_159_224 ();
 FILLCELL_X32 FILLCELL_159_256 ();
 FILLCELL_X32 FILLCELL_159_288 ();
 FILLCELL_X32 FILLCELL_159_320 ();
 FILLCELL_X32 FILLCELL_159_352 ();
 FILLCELL_X32 FILLCELL_159_384 ();
 FILLCELL_X32 FILLCELL_159_416 ();
 FILLCELL_X32 FILLCELL_159_448 ();
 FILLCELL_X32 FILLCELL_159_480 ();
 FILLCELL_X32 FILLCELL_159_512 ();
 FILLCELL_X32 FILLCELL_159_544 ();
 FILLCELL_X32 FILLCELL_159_576 ();
 FILLCELL_X32 FILLCELL_159_608 ();
 FILLCELL_X32 FILLCELL_159_640 ();
 FILLCELL_X32 FILLCELL_159_672 ();
 FILLCELL_X32 FILLCELL_159_704 ();
 FILLCELL_X32 FILLCELL_159_736 ();
 FILLCELL_X32 FILLCELL_159_768 ();
 FILLCELL_X32 FILLCELL_159_800 ();
 FILLCELL_X32 FILLCELL_159_832 ();
 FILLCELL_X32 FILLCELL_159_864 ();
 FILLCELL_X32 FILLCELL_159_896 ();
 FILLCELL_X32 FILLCELL_159_928 ();
 FILLCELL_X32 FILLCELL_159_960 ();
 FILLCELL_X32 FILLCELL_159_992 ();
 FILLCELL_X32 FILLCELL_159_1024 ();
 FILLCELL_X32 FILLCELL_159_1056 ();
 FILLCELL_X32 FILLCELL_159_1088 ();
 FILLCELL_X32 FILLCELL_159_1120 ();
 FILLCELL_X32 FILLCELL_159_1152 ();
 FILLCELL_X32 FILLCELL_159_1184 ();
 FILLCELL_X32 FILLCELL_159_1216 ();
 FILLCELL_X32 FILLCELL_159_1248 ();
 FILLCELL_X32 FILLCELL_159_1280 ();
 FILLCELL_X32 FILLCELL_159_1312 ();
 FILLCELL_X32 FILLCELL_159_1344 ();
 FILLCELL_X32 FILLCELL_159_1376 ();
 FILLCELL_X32 FILLCELL_159_1408 ();
 FILLCELL_X32 FILLCELL_159_1440 ();
 FILLCELL_X32 FILLCELL_159_1472 ();
 FILLCELL_X32 FILLCELL_159_1504 ();
 FILLCELL_X32 FILLCELL_159_1536 ();
 FILLCELL_X32 FILLCELL_159_1568 ();
 FILLCELL_X32 FILLCELL_159_1600 ();
 FILLCELL_X32 FILLCELL_159_1632 ();
 FILLCELL_X32 FILLCELL_159_1664 ();
 FILLCELL_X32 FILLCELL_159_1696 ();
 FILLCELL_X32 FILLCELL_159_1728 ();
 FILLCELL_X32 FILLCELL_159_1760 ();
 FILLCELL_X32 FILLCELL_159_1792 ();
 FILLCELL_X32 FILLCELL_159_1824 ();
 FILLCELL_X32 FILLCELL_159_1856 ();
 FILLCELL_X8 FILLCELL_159_1888 ();
 FILLCELL_X1 FILLCELL_159_1896 ();
 FILLCELL_X32 FILLCELL_160_0 ();
 FILLCELL_X32 FILLCELL_160_32 ();
 FILLCELL_X32 FILLCELL_160_64 ();
 FILLCELL_X32 FILLCELL_160_96 ();
 FILLCELL_X32 FILLCELL_160_128 ();
 FILLCELL_X4 FILLCELL_160_160 ();
 FILLCELL_X32 FILLCELL_160_167 ();
 FILLCELL_X32 FILLCELL_160_199 ();
 FILLCELL_X32 FILLCELL_160_231 ();
 FILLCELL_X32 FILLCELL_160_263 ();
 FILLCELL_X32 FILLCELL_160_295 ();
 FILLCELL_X32 FILLCELL_160_327 ();
 FILLCELL_X32 FILLCELL_160_359 ();
 FILLCELL_X32 FILLCELL_160_391 ();
 FILLCELL_X32 FILLCELL_160_423 ();
 FILLCELL_X32 FILLCELL_160_455 ();
 FILLCELL_X32 FILLCELL_160_487 ();
 FILLCELL_X32 FILLCELL_160_519 ();
 FILLCELL_X32 FILLCELL_160_551 ();
 FILLCELL_X32 FILLCELL_160_583 ();
 FILLCELL_X32 FILLCELL_160_615 ();
 FILLCELL_X32 FILLCELL_160_647 ();
 FILLCELL_X32 FILLCELL_160_679 ();
 FILLCELL_X16 FILLCELL_160_711 ();
 FILLCELL_X32 FILLCELL_160_732 ();
 FILLCELL_X32 FILLCELL_160_764 ();
 FILLCELL_X16 FILLCELL_160_796 ();
 FILLCELL_X8 FILLCELL_160_812 ();
 FILLCELL_X4 FILLCELL_160_820 ();
 FILLCELL_X2 FILLCELL_160_824 ();
 FILLCELL_X1 FILLCELL_160_826 ();
 FILLCELL_X32 FILLCELL_160_830 ();
 FILLCELL_X32 FILLCELL_160_862 ();
 FILLCELL_X32 FILLCELL_160_894 ();
 FILLCELL_X32 FILLCELL_160_926 ();
 FILLCELL_X32 FILLCELL_160_958 ();
 FILLCELL_X32 FILLCELL_160_990 ();
 FILLCELL_X32 FILLCELL_160_1022 ();
 FILLCELL_X32 FILLCELL_160_1054 ();
 FILLCELL_X32 FILLCELL_160_1086 ();
 FILLCELL_X32 FILLCELL_160_1118 ();
 FILLCELL_X32 FILLCELL_160_1150 ();
 FILLCELL_X32 FILLCELL_160_1182 ();
 FILLCELL_X32 FILLCELL_160_1214 ();
 FILLCELL_X32 FILLCELL_160_1246 ();
 FILLCELL_X32 FILLCELL_160_1278 ();
 FILLCELL_X32 FILLCELL_160_1310 ();
 FILLCELL_X32 FILLCELL_160_1342 ();
 FILLCELL_X32 FILLCELL_160_1374 ();
 FILLCELL_X32 FILLCELL_160_1406 ();
 FILLCELL_X32 FILLCELL_160_1438 ();
 FILLCELL_X32 FILLCELL_160_1470 ();
 FILLCELL_X32 FILLCELL_160_1502 ();
 FILLCELL_X32 FILLCELL_160_1534 ();
 FILLCELL_X32 FILLCELL_160_1566 ();
 FILLCELL_X32 FILLCELL_160_1598 ();
 FILLCELL_X32 FILLCELL_160_1630 ();
 FILLCELL_X32 FILLCELL_160_1662 ();
 FILLCELL_X32 FILLCELL_160_1694 ();
 FILLCELL_X32 FILLCELL_160_1726 ();
 FILLCELL_X32 FILLCELL_160_1758 ();
 FILLCELL_X32 FILLCELL_160_1790 ();
 FILLCELL_X32 FILLCELL_160_1822 ();
 FILLCELL_X32 FILLCELL_160_1854 ();
 FILLCELL_X8 FILLCELL_160_1886 ();
 FILLCELL_X2 FILLCELL_160_1894 ();
 FILLCELL_X1 FILLCELL_160_1896 ();
 FILLCELL_X32 FILLCELL_161_0 ();
 FILLCELL_X32 FILLCELL_161_32 ();
 FILLCELL_X4 FILLCELL_161_64 ();
 FILLCELL_X32 FILLCELL_161_85 ();
 FILLCELL_X32 FILLCELL_161_117 ();
 FILLCELL_X32 FILLCELL_161_149 ();
 FILLCELL_X32 FILLCELL_161_181 ();
 FILLCELL_X32 FILLCELL_161_213 ();
 FILLCELL_X32 FILLCELL_161_245 ();
 FILLCELL_X32 FILLCELL_161_277 ();
 FILLCELL_X32 FILLCELL_161_309 ();
 FILLCELL_X32 FILLCELL_161_341 ();
 FILLCELL_X32 FILLCELL_161_373 ();
 FILLCELL_X32 FILLCELL_161_405 ();
 FILLCELL_X32 FILLCELL_161_437 ();
 FILLCELL_X32 FILLCELL_161_469 ();
 FILLCELL_X32 FILLCELL_161_501 ();
 FILLCELL_X32 FILLCELL_161_533 ();
 FILLCELL_X32 FILLCELL_161_565 ();
 FILLCELL_X32 FILLCELL_161_597 ();
 FILLCELL_X32 FILLCELL_161_629 ();
 FILLCELL_X32 FILLCELL_161_661 ();
 FILLCELL_X32 FILLCELL_161_693 ();
 FILLCELL_X8 FILLCELL_161_725 ();
 FILLCELL_X2 FILLCELL_161_733 ();
 FILLCELL_X1 FILLCELL_161_735 ();
 FILLCELL_X32 FILLCELL_161_741 ();
 FILLCELL_X32 FILLCELL_161_773 ();
 FILLCELL_X32 FILLCELL_161_805 ();
 FILLCELL_X32 FILLCELL_161_837 ();
 FILLCELL_X32 FILLCELL_161_869 ();
 FILLCELL_X32 FILLCELL_161_901 ();
 FILLCELL_X32 FILLCELL_161_933 ();
 FILLCELL_X8 FILLCELL_161_965 ();
 FILLCELL_X4 FILLCELL_161_973 ();
 FILLCELL_X2 FILLCELL_161_977 ();
 FILLCELL_X1 FILLCELL_161_979 ();
 FILLCELL_X32 FILLCELL_161_985 ();
 FILLCELL_X32 FILLCELL_161_1017 ();
 FILLCELL_X32 FILLCELL_161_1049 ();
 FILLCELL_X2 FILLCELL_161_1081 ();
 FILLCELL_X32 FILLCELL_161_1086 ();
 FILLCELL_X32 FILLCELL_161_1118 ();
 FILLCELL_X32 FILLCELL_161_1150 ();
 FILLCELL_X32 FILLCELL_161_1182 ();
 FILLCELL_X32 FILLCELL_161_1214 ();
 FILLCELL_X32 FILLCELL_161_1246 ();
 FILLCELL_X32 FILLCELL_161_1278 ();
 FILLCELL_X32 FILLCELL_161_1310 ();
 FILLCELL_X32 FILLCELL_161_1342 ();
 FILLCELL_X32 FILLCELL_161_1374 ();
 FILLCELL_X32 FILLCELL_161_1406 ();
 FILLCELL_X32 FILLCELL_161_1438 ();
 FILLCELL_X32 FILLCELL_161_1470 ();
 FILLCELL_X32 FILLCELL_161_1502 ();
 FILLCELL_X32 FILLCELL_161_1534 ();
 FILLCELL_X32 FILLCELL_161_1566 ();
 FILLCELL_X32 FILLCELL_161_1598 ();
 FILLCELL_X32 FILLCELL_161_1630 ();
 FILLCELL_X32 FILLCELL_161_1662 ();
 FILLCELL_X32 FILLCELL_161_1694 ();
 FILLCELL_X32 FILLCELL_161_1726 ();
 FILLCELL_X32 FILLCELL_161_1758 ();
 FILLCELL_X32 FILLCELL_161_1790 ();
 FILLCELL_X32 FILLCELL_161_1822 ();
 FILLCELL_X32 FILLCELL_161_1854 ();
 FILLCELL_X8 FILLCELL_161_1886 ();
 FILLCELL_X2 FILLCELL_161_1894 ();
 FILLCELL_X1 FILLCELL_161_1896 ();
 FILLCELL_X32 FILLCELL_162_0 ();
 FILLCELL_X32 FILLCELL_162_32 ();
 FILLCELL_X32 FILLCELL_162_64 ();
 FILLCELL_X32 FILLCELL_162_96 ();
 FILLCELL_X4 FILLCELL_162_128 ();
 FILLCELL_X32 FILLCELL_162_135 ();
 FILLCELL_X32 FILLCELL_162_167 ();
 FILLCELL_X32 FILLCELL_162_199 ();
 FILLCELL_X32 FILLCELL_162_231 ();
 FILLCELL_X32 FILLCELL_162_263 ();
 FILLCELL_X32 FILLCELL_162_295 ();
 FILLCELL_X32 FILLCELL_162_327 ();
 FILLCELL_X32 FILLCELL_162_359 ();
 FILLCELL_X32 FILLCELL_162_391 ();
 FILLCELL_X32 FILLCELL_162_423 ();
 FILLCELL_X32 FILLCELL_162_455 ();
 FILLCELL_X32 FILLCELL_162_487 ();
 FILLCELL_X32 FILLCELL_162_519 ();
 FILLCELL_X32 FILLCELL_162_551 ();
 FILLCELL_X32 FILLCELL_162_583 ();
 FILLCELL_X32 FILLCELL_162_615 ();
 FILLCELL_X32 FILLCELL_162_647 ();
 FILLCELL_X32 FILLCELL_162_679 ();
 FILLCELL_X32 FILLCELL_162_711 ();
 FILLCELL_X32 FILLCELL_162_743 ();
 FILLCELL_X32 FILLCELL_162_775 ();
 FILLCELL_X32 FILLCELL_162_807 ();
 FILLCELL_X32 FILLCELL_162_839 ();
 FILLCELL_X32 FILLCELL_162_871 ();
 FILLCELL_X32 FILLCELL_162_903 ();
 FILLCELL_X32 FILLCELL_162_935 ();
 FILLCELL_X16 FILLCELL_162_967 ();
 FILLCELL_X8 FILLCELL_162_983 ();
 FILLCELL_X2 FILLCELL_162_991 ();
 FILLCELL_X32 FILLCELL_162_1002 ();
 FILLCELL_X32 FILLCELL_162_1034 ();
 FILLCELL_X32 FILLCELL_162_1066 ();
 FILLCELL_X32 FILLCELL_162_1098 ();
 FILLCELL_X32 FILLCELL_162_1130 ();
 FILLCELL_X32 FILLCELL_162_1162 ();
 FILLCELL_X32 FILLCELL_162_1194 ();
 FILLCELL_X32 FILLCELL_162_1226 ();
 FILLCELL_X32 FILLCELL_162_1258 ();
 FILLCELL_X32 FILLCELL_162_1290 ();
 FILLCELL_X32 FILLCELL_162_1322 ();
 FILLCELL_X32 FILLCELL_162_1354 ();
 FILLCELL_X32 FILLCELL_162_1386 ();
 FILLCELL_X32 FILLCELL_162_1418 ();
 FILLCELL_X32 FILLCELL_162_1450 ();
 FILLCELL_X32 FILLCELL_162_1482 ();
 FILLCELL_X32 FILLCELL_162_1514 ();
 FILLCELL_X32 FILLCELL_162_1546 ();
 FILLCELL_X32 FILLCELL_162_1578 ();
 FILLCELL_X32 FILLCELL_162_1610 ();
 FILLCELL_X32 FILLCELL_162_1642 ();
 FILLCELL_X32 FILLCELL_162_1674 ();
 FILLCELL_X32 FILLCELL_162_1706 ();
 FILLCELL_X32 FILLCELL_162_1738 ();
 FILLCELL_X32 FILLCELL_162_1770 ();
 FILLCELL_X32 FILLCELL_162_1802 ();
 FILLCELL_X32 FILLCELL_162_1834 ();
 FILLCELL_X16 FILLCELL_162_1866 ();
 FILLCELL_X8 FILLCELL_162_1882 ();
 FILLCELL_X4 FILLCELL_162_1890 ();
 FILLCELL_X2 FILLCELL_162_1894 ();
 FILLCELL_X1 FILLCELL_162_1896 ();
 FILLCELL_X32 FILLCELL_163_0 ();
 FILLCELL_X32 FILLCELL_163_32 ();
 FILLCELL_X32 FILLCELL_163_64 ();
 FILLCELL_X32 FILLCELL_163_96 ();
 FILLCELL_X32 FILLCELL_163_128 ();
 FILLCELL_X32 FILLCELL_163_160 ();
 FILLCELL_X32 FILLCELL_163_192 ();
 FILLCELL_X32 FILLCELL_163_224 ();
 FILLCELL_X32 FILLCELL_163_256 ();
 FILLCELL_X16 FILLCELL_163_288 ();
 FILLCELL_X2 FILLCELL_163_304 ();
 FILLCELL_X1 FILLCELL_163_306 ();
 FILLCELL_X32 FILLCELL_163_310 ();
 FILLCELL_X32 FILLCELL_163_342 ();
 FILLCELL_X32 FILLCELL_163_374 ();
 FILLCELL_X32 FILLCELL_163_406 ();
 FILLCELL_X32 FILLCELL_163_438 ();
 FILLCELL_X32 FILLCELL_163_470 ();
 FILLCELL_X32 FILLCELL_163_502 ();
 FILLCELL_X32 FILLCELL_163_534 ();
 FILLCELL_X32 FILLCELL_163_566 ();
 FILLCELL_X32 FILLCELL_163_598 ();
 FILLCELL_X32 FILLCELL_163_630 ();
 FILLCELL_X16 FILLCELL_163_662 ();
 FILLCELL_X2 FILLCELL_163_678 ();
 FILLCELL_X1 FILLCELL_163_680 ();
 FILLCELL_X32 FILLCELL_163_683 ();
 FILLCELL_X32 FILLCELL_163_715 ();
 FILLCELL_X32 FILLCELL_163_747 ();
 FILLCELL_X32 FILLCELL_163_779 ();
 FILLCELL_X32 FILLCELL_163_811 ();
 FILLCELL_X32 FILLCELL_163_843 ();
 FILLCELL_X32 FILLCELL_163_875 ();
 FILLCELL_X32 FILLCELL_163_907 ();
 FILLCELL_X32 FILLCELL_163_939 ();
 FILLCELL_X32 FILLCELL_163_971 ();
 FILLCELL_X32 FILLCELL_163_1003 ();
 FILLCELL_X32 FILLCELL_163_1035 ();
 FILLCELL_X32 FILLCELL_163_1067 ();
 FILLCELL_X32 FILLCELL_163_1099 ();
 FILLCELL_X32 FILLCELL_163_1131 ();
 FILLCELL_X32 FILLCELL_163_1163 ();
 FILLCELL_X32 FILLCELL_163_1195 ();
 FILLCELL_X32 FILLCELL_163_1227 ();
 FILLCELL_X32 FILLCELL_163_1259 ();
 FILLCELL_X32 FILLCELL_163_1291 ();
 FILLCELL_X32 FILLCELL_163_1323 ();
 FILLCELL_X32 FILLCELL_163_1355 ();
 FILLCELL_X32 FILLCELL_163_1387 ();
 FILLCELL_X32 FILLCELL_163_1419 ();
 FILLCELL_X32 FILLCELL_163_1451 ();
 FILLCELL_X32 FILLCELL_163_1483 ();
 FILLCELL_X32 FILLCELL_163_1515 ();
 FILLCELL_X32 FILLCELL_163_1547 ();
 FILLCELL_X32 FILLCELL_163_1579 ();
 FILLCELL_X32 FILLCELL_163_1611 ();
 FILLCELL_X32 FILLCELL_163_1643 ();
 FILLCELL_X32 FILLCELL_163_1675 ();
 FILLCELL_X32 FILLCELL_163_1707 ();
 FILLCELL_X32 FILLCELL_163_1739 ();
 FILLCELL_X32 FILLCELL_163_1771 ();
 FILLCELL_X32 FILLCELL_163_1803 ();
 FILLCELL_X32 FILLCELL_163_1835 ();
 FILLCELL_X16 FILLCELL_163_1867 ();
 FILLCELL_X8 FILLCELL_163_1883 ();
 FILLCELL_X4 FILLCELL_163_1891 ();
 FILLCELL_X2 FILLCELL_163_1895 ();
 FILLCELL_X32 FILLCELL_164_0 ();
 FILLCELL_X32 FILLCELL_164_32 ();
 FILLCELL_X32 FILLCELL_164_64 ();
 FILLCELL_X32 FILLCELL_164_96 ();
 FILLCELL_X32 FILLCELL_164_128 ();
 FILLCELL_X32 FILLCELL_164_160 ();
 FILLCELL_X32 FILLCELL_164_192 ();
 FILLCELL_X32 FILLCELL_164_224 ();
 FILLCELL_X32 FILLCELL_164_256 ();
 FILLCELL_X32 FILLCELL_164_288 ();
 FILLCELL_X32 FILLCELL_164_320 ();
 FILLCELL_X32 FILLCELL_164_352 ();
 FILLCELL_X8 FILLCELL_164_384 ();
 FILLCELL_X4 FILLCELL_164_392 ();
 FILLCELL_X32 FILLCELL_164_405 ();
 FILLCELL_X32 FILLCELL_164_437 ();
 FILLCELL_X16 FILLCELL_164_469 ();
 FILLCELL_X8 FILLCELL_164_485 ();
 FILLCELL_X32 FILLCELL_164_495 ();
 FILLCELL_X16 FILLCELL_164_527 ();
 FILLCELL_X8 FILLCELL_164_543 ();
 FILLCELL_X4 FILLCELL_164_551 ();
 FILLCELL_X1 FILLCELL_164_555 ();
 FILLCELL_X4 FILLCELL_164_559 ();
 FILLCELL_X8 FILLCELL_164_569 ();
 FILLCELL_X2 FILLCELL_164_577 ();
 FILLCELL_X1 FILLCELL_164_579 ();
 FILLCELL_X8 FILLCELL_164_584 ();
 FILLCELL_X4 FILLCELL_164_592 ();
 FILLCELL_X32 FILLCELL_164_605 ();
 FILLCELL_X32 FILLCELL_164_637 ();
 FILLCELL_X32 FILLCELL_164_669 ();
 FILLCELL_X32 FILLCELL_164_701 ();
 FILLCELL_X32 FILLCELL_164_733 ();
 FILLCELL_X32 FILLCELL_164_765 ();
 FILLCELL_X16 FILLCELL_164_797 ();
 FILLCELL_X4 FILLCELL_164_813 ();
 FILLCELL_X2 FILLCELL_164_817 ();
 FILLCELL_X32 FILLCELL_164_822 ();
 FILLCELL_X32 FILLCELL_164_854 ();
 FILLCELL_X32 FILLCELL_164_886 ();
 FILLCELL_X32 FILLCELL_164_918 ();
 FILLCELL_X32 FILLCELL_164_950 ();
 FILLCELL_X32 FILLCELL_164_982 ();
 FILLCELL_X32 FILLCELL_164_1014 ();
 FILLCELL_X32 FILLCELL_164_1046 ();
 FILLCELL_X32 FILLCELL_164_1078 ();
 FILLCELL_X32 FILLCELL_164_1110 ();
 FILLCELL_X32 FILLCELL_164_1142 ();
 FILLCELL_X32 FILLCELL_164_1174 ();
 FILLCELL_X32 FILLCELL_164_1206 ();
 FILLCELL_X32 FILLCELL_164_1238 ();
 FILLCELL_X32 FILLCELL_164_1270 ();
 FILLCELL_X32 FILLCELL_164_1302 ();
 FILLCELL_X32 FILLCELL_164_1334 ();
 FILLCELL_X32 FILLCELL_164_1366 ();
 FILLCELL_X32 FILLCELL_164_1398 ();
 FILLCELL_X32 FILLCELL_164_1430 ();
 FILLCELL_X32 FILLCELL_164_1462 ();
 FILLCELL_X32 FILLCELL_164_1494 ();
 FILLCELL_X32 FILLCELL_164_1526 ();
 FILLCELL_X32 FILLCELL_164_1558 ();
 FILLCELL_X32 FILLCELL_164_1590 ();
 FILLCELL_X32 FILLCELL_164_1622 ();
 FILLCELL_X32 FILLCELL_164_1654 ();
 FILLCELL_X32 FILLCELL_164_1686 ();
 FILLCELL_X32 FILLCELL_164_1718 ();
 FILLCELL_X32 FILLCELL_164_1750 ();
 FILLCELL_X32 FILLCELL_164_1782 ();
 FILLCELL_X32 FILLCELL_164_1814 ();
 FILLCELL_X32 FILLCELL_164_1846 ();
 FILLCELL_X16 FILLCELL_164_1878 ();
 FILLCELL_X2 FILLCELL_164_1894 ();
 FILLCELL_X1 FILLCELL_164_1896 ();
 FILLCELL_X32 FILLCELL_165_0 ();
 FILLCELL_X32 FILLCELL_165_32 ();
 FILLCELL_X32 FILLCELL_165_64 ();
 FILLCELL_X32 FILLCELL_165_96 ();
 FILLCELL_X32 FILLCELL_165_128 ();
 FILLCELL_X32 FILLCELL_165_160 ();
 FILLCELL_X32 FILLCELL_165_192 ();
 FILLCELL_X32 FILLCELL_165_224 ();
 FILLCELL_X32 FILLCELL_165_256 ();
 FILLCELL_X32 FILLCELL_165_288 ();
 FILLCELL_X32 FILLCELL_165_320 ();
 FILLCELL_X32 FILLCELL_165_352 ();
 FILLCELL_X16 FILLCELL_165_384 ();
 FILLCELL_X8 FILLCELL_165_400 ();
 FILLCELL_X4 FILLCELL_165_408 ();
 FILLCELL_X2 FILLCELL_165_412 ();
 FILLCELL_X32 FILLCELL_165_418 ();
 FILLCELL_X32 FILLCELL_165_450 ();
 FILLCELL_X32 FILLCELL_165_482 ();
 FILLCELL_X32 FILLCELL_165_514 ();
 FILLCELL_X32 FILLCELL_165_546 ();
 FILLCELL_X32 FILLCELL_165_578 ();
 FILLCELL_X32 FILLCELL_165_610 ();
 FILLCELL_X32 FILLCELL_165_642 ();
 FILLCELL_X32 FILLCELL_165_674 ();
 FILLCELL_X32 FILLCELL_165_706 ();
 FILLCELL_X32 FILLCELL_165_738 ();
 FILLCELL_X32 FILLCELL_165_770 ();
 FILLCELL_X32 FILLCELL_165_802 ();
 FILLCELL_X32 FILLCELL_165_834 ();
 FILLCELL_X32 FILLCELL_165_866 ();
 FILLCELL_X16 FILLCELL_165_898 ();
 FILLCELL_X1 FILLCELL_165_914 ();
 FILLCELL_X32 FILLCELL_165_918 ();
 FILLCELL_X32 FILLCELL_165_950 ();
 FILLCELL_X32 FILLCELL_165_982 ();
 FILLCELL_X32 FILLCELL_165_1014 ();
 FILLCELL_X32 FILLCELL_165_1046 ();
 FILLCELL_X32 FILLCELL_165_1078 ();
 FILLCELL_X32 FILLCELL_165_1110 ();
 FILLCELL_X32 FILLCELL_165_1142 ();
 FILLCELL_X32 FILLCELL_165_1174 ();
 FILLCELL_X32 FILLCELL_165_1206 ();
 FILLCELL_X32 FILLCELL_165_1238 ();
 FILLCELL_X32 FILLCELL_165_1270 ();
 FILLCELL_X32 FILLCELL_165_1302 ();
 FILLCELL_X32 FILLCELL_165_1334 ();
 FILLCELL_X32 FILLCELL_165_1366 ();
 FILLCELL_X32 FILLCELL_165_1398 ();
 FILLCELL_X32 FILLCELL_165_1430 ();
 FILLCELL_X32 FILLCELL_165_1462 ();
 FILLCELL_X32 FILLCELL_165_1494 ();
 FILLCELL_X32 FILLCELL_165_1526 ();
 FILLCELL_X32 FILLCELL_165_1558 ();
 FILLCELL_X32 FILLCELL_165_1590 ();
 FILLCELL_X32 FILLCELL_165_1622 ();
 FILLCELL_X32 FILLCELL_165_1654 ();
 FILLCELL_X32 FILLCELL_165_1686 ();
 FILLCELL_X32 FILLCELL_165_1718 ();
 FILLCELL_X32 FILLCELL_165_1750 ();
 FILLCELL_X32 FILLCELL_165_1782 ();
 FILLCELL_X32 FILLCELL_165_1814 ();
 FILLCELL_X32 FILLCELL_165_1846 ();
 FILLCELL_X16 FILLCELL_165_1878 ();
 FILLCELL_X2 FILLCELL_165_1894 ();
 FILLCELL_X1 FILLCELL_165_1896 ();
 FILLCELL_X32 FILLCELL_166_0 ();
 FILLCELL_X32 FILLCELL_166_32 ();
 FILLCELL_X32 FILLCELL_166_64 ();
 FILLCELL_X32 FILLCELL_166_96 ();
 FILLCELL_X32 FILLCELL_166_128 ();
 FILLCELL_X32 FILLCELL_166_160 ();
 FILLCELL_X16 FILLCELL_166_192 ();
 FILLCELL_X32 FILLCELL_166_215 ();
 FILLCELL_X32 FILLCELL_166_247 ();
 FILLCELL_X32 FILLCELL_166_279 ();
 FILLCELL_X32 FILLCELL_166_311 ();
 FILLCELL_X32 FILLCELL_166_343 ();
 FILLCELL_X32 FILLCELL_166_375 ();
 FILLCELL_X32 FILLCELL_166_407 ();
 FILLCELL_X32 FILLCELL_166_439 ();
 FILLCELL_X1 FILLCELL_166_471 ();
 FILLCELL_X32 FILLCELL_166_485 ();
 FILLCELL_X32 FILLCELL_166_517 ();
 FILLCELL_X32 FILLCELL_166_549 ();
 FILLCELL_X32 FILLCELL_166_581 ();
 FILLCELL_X32 FILLCELL_166_613 ();
 FILLCELL_X16 FILLCELL_166_645 ();
 FILLCELL_X8 FILLCELL_166_661 ();
 FILLCELL_X2 FILLCELL_166_669 ();
 FILLCELL_X32 FILLCELL_166_678 ();
 FILLCELL_X16 FILLCELL_166_710 ();
 FILLCELL_X8 FILLCELL_166_726 ();
 FILLCELL_X4 FILLCELL_166_734 ();
 FILLCELL_X32 FILLCELL_166_740 ();
 FILLCELL_X32 FILLCELL_166_772 ();
 FILLCELL_X16 FILLCELL_166_804 ();
 FILLCELL_X4 FILLCELL_166_820 ();
 FILLCELL_X2 FILLCELL_166_824 ();
 FILLCELL_X1 FILLCELL_166_826 ();
 FILLCELL_X4 FILLCELL_166_830 ();
 FILLCELL_X32 FILLCELL_166_838 ();
 FILLCELL_X32 FILLCELL_166_870 ();
 FILLCELL_X32 FILLCELL_166_902 ();
 FILLCELL_X32 FILLCELL_166_934 ();
 FILLCELL_X32 FILLCELL_166_966 ();
 FILLCELL_X32 FILLCELL_166_998 ();
 FILLCELL_X32 FILLCELL_166_1030 ();
 FILLCELL_X32 FILLCELL_166_1062 ();
 FILLCELL_X32 FILLCELL_166_1094 ();
 FILLCELL_X32 FILLCELL_166_1126 ();
 FILLCELL_X32 FILLCELL_166_1158 ();
 FILLCELL_X32 FILLCELL_166_1190 ();
 FILLCELL_X32 FILLCELL_166_1222 ();
 FILLCELL_X32 FILLCELL_166_1254 ();
 FILLCELL_X32 FILLCELL_166_1286 ();
 FILLCELL_X32 FILLCELL_166_1318 ();
 FILLCELL_X32 FILLCELL_166_1350 ();
 FILLCELL_X32 FILLCELL_166_1382 ();
 FILLCELL_X32 FILLCELL_166_1414 ();
 FILLCELL_X32 FILLCELL_166_1446 ();
 FILLCELL_X32 FILLCELL_166_1478 ();
 FILLCELL_X32 FILLCELL_166_1510 ();
 FILLCELL_X32 FILLCELL_166_1542 ();
 FILLCELL_X32 FILLCELL_166_1574 ();
 FILLCELL_X32 FILLCELL_166_1606 ();
 FILLCELL_X32 FILLCELL_166_1638 ();
 FILLCELL_X32 FILLCELL_166_1670 ();
 FILLCELL_X32 FILLCELL_166_1702 ();
 FILLCELL_X32 FILLCELL_166_1734 ();
 FILLCELL_X32 FILLCELL_166_1766 ();
 FILLCELL_X32 FILLCELL_166_1798 ();
 FILLCELL_X32 FILLCELL_166_1830 ();
 FILLCELL_X32 FILLCELL_166_1862 ();
 FILLCELL_X2 FILLCELL_166_1894 ();
 FILLCELL_X1 FILLCELL_166_1896 ();
 FILLCELL_X32 FILLCELL_167_0 ();
 FILLCELL_X32 FILLCELL_167_32 ();
 FILLCELL_X32 FILLCELL_167_64 ();
 FILLCELL_X32 FILLCELL_167_96 ();
 FILLCELL_X32 FILLCELL_167_128 ();
 FILLCELL_X32 FILLCELL_167_160 ();
 FILLCELL_X32 FILLCELL_167_192 ();
 FILLCELL_X32 FILLCELL_167_224 ();
 FILLCELL_X4 FILLCELL_167_256 ();
 FILLCELL_X2 FILLCELL_167_260 ();
 FILLCELL_X1 FILLCELL_167_262 ();
 FILLCELL_X32 FILLCELL_167_280 ();
 FILLCELL_X32 FILLCELL_167_312 ();
 FILLCELL_X32 FILLCELL_167_344 ();
 FILLCELL_X32 FILLCELL_167_376 ();
 FILLCELL_X32 FILLCELL_167_408 ();
 FILLCELL_X32 FILLCELL_167_440 ();
 FILLCELL_X8 FILLCELL_167_472 ();
 FILLCELL_X32 FILLCELL_167_482 ();
 FILLCELL_X32 FILLCELL_167_514 ();
 FILLCELL_X32 FILLCELL_167_546 ();
 FILLCELL_X32 FILLCELL_167_578 ();
 FILLCELL_X32 FILLCELL_167_610 ();
 FILLCELL_X16 FILLCELL_167_642 ();
 FILLCELL_X4 FILLCELL_167_658 ();
 FILLCELL_X2 FILLCELL_167_662 ();
 FILLCELL_X32 FILLCELL_167_666 ();
 FILLCELL_X32 FILLCELL_167_698 ();
 FILLCELL_X32 FILLCELL_167_730 ();
 FILLCELL_X32 FILLCELL_167_762 ();
 FILLCELL_X32 FILLCELL_167_794 ();
 FILLCELL_X8 FILLCELL_167_826 ();
 FILLCELL_X32 FILLCELL_167_836 ();
 FILLCELL_X32 FILLCELL_167_868 ();
 FILLCELL_X32 FILLCELL_167_900 ();
 FILLCELL_X32 FILLCELL_167_932 ();
 FILLCELL_X32 FILLCELL_167_964 ();
 FILLCELL_X32 FILLCELL_167_996 ();
 FILLCELL_X32 FILLCELL_167_1028 ();
 FILLCELL_X32 FILLCELL_167_1060 ();
 FILLCELL_X32 FILLCELL_167_1092 ();
 FILLCELL_X4 FILLCELL_167_1124 ();
 FILLCELL_X2 FILLCELL_167_1128 ();
 FILLCELL_X32 FILLCELL_167_1143 ();
 FILLCELL_X32 FILLCELL_167_1175 ();
 FILLCELL_X32 FILLCELL_167_1207 ();
 FILLCELL_X32 FILLCELL_167_1239 ();
 FILLCELL_X32 FILLCELL_167_1271 ();
 FILLCELL_X32 FILLCELL_167_1303 ();
 FILLCELL_X32 FILLCELL_167_1335 ();
 FILLCELL_X32 FILLCELL_167_1367 ();
 FILLCELL_X32 FILLCELL_167_1399 ();
 FILLCELL_X32 FILLCELL_167_1431 ();
 FILLCELL_X32 FILLCELL_167_1463 ();
 FILLCELL_X32 FILLCELL_167_1495 ();
 FILLCELL_X32 FILLCELL_167_1527 ();
 FILLCELL_X32 FILLCELL_167_1559 ();
 FILLCELL_X32 FILLCELL_167_1591 ();
 FILLCELL_X32 FILLCELL_167_1623 ();
 FILLCELL_X32 FILLCELL_167_1655 ();
 FILLCELL_X32 FILLCELL_167_1687 ();
 FILLCELL_X32 FILLCELL_167_1719 ();
 FILLCELL_X32 FILLCELL_167_1751 ();
 FILLCELL_X32 FILLCELL_167_1783 ();
 FILLCELL_X32 FILLCELL_167_1815 ();
 FILLCELL_X32 FILLCELL_167_1847 ();
 FILLCELL_X16 FILLCELL_167_1879 ();
 FILLCELL_X2 FILLCELL_167_1895 ();
 FILLCELL_X32 FILLCELL_168_0 ();
 FILLCELL_X32 FILLCELL_168_32 ();
 FILLCELL_X32 FILLCELL_168_64 ();
 FILLCELL_X32 FILLCELL_168_96 ();
 FILLCELL_X32 FILLCELL_168_128 ();
 FILLCELL_X32 FILLCELL_168_160 ();
 FILLCELL_X32 FILLCELL_168_192 ();
 FILLCELL_X32 FILLCELL_168_224 ();
 FILLCELL_X32 FILLCELL_168_256 ();
 FILLCELL_X32 FILLCELL_168_288 ();
 FILLCELL_X32 FILLCELL_168_320 ();
 FILLCELL_X32 FILLCELL_168_352 ();
 FILLCELL_X8 FILLCELL_168_384 ();
 FILLCELL_X1 FILLCELL_168_392 ();
 FILLCELL_X32 FILLCELL_168_396 ();
 FILLCELL_X2 FILLCELL_168_428 ();
 FILLCELL_X32 FILLCELL_168_435 ();
 FILLCELL_X32 FILLCELL_168_467 ();
 FILLCELL_X32 FILLCELL_168_499 ();
 FILLCELL_X32 FILLCELL_168_531 ();
 FILLCELL_X32 FILLCELL_168_563 ();
 FILLCELL_X32 FILLCELL_168_595 ();
 FILLCELL_X32 FILLCELL_168_627 ();
 FILLCELL_X32 FILLCELL_168_659 ();
 FILLCELL_X32 FILLCELL_168_691 ();
 FILLCELL_X32 FILLCELL_168_723 ();
 FILLCELL_X32 FILLCELL_168_755 ();
 FILLCELL_X32 FILLCELL_168_787 ();
 FILLCELL_X16 FILLCELL_168_819 ();
 FILLCELL_X8 FILLCELL_168_835 ();
 FILLCELL_X2 FILLCELL_168_843 ();
 FILLCELL_X1 FILLCELL_168_845 ();
 FILLCELL_X32 FILLCELL_168_849 ();
 FILLCELL_X16 FILLCELL_168_881 ();
 FILLCELL_X4 FILLCELL_168_897 ();
 FILLCELL_X1 FILLCELL_168_901 ();
 FILLCELL_X32 FILLCELL_168_906 ();
 FILLCELL_X32 FILLCELL_168_938 ();
 FILLCELL_X8 FILLCELL_168_970 ();
 FILLCELL_X2 FILLCELL_168_978 ();
 FILLCELL_X1 FILLCELL_168_980 ();
 FILLCELL_X32 FILLCELL_168_988 ();
 FILLCELL_X32 FILLCELL_168_1020 ();
 FILLCELL_X32 FILLCELL_168_1052 ();
 FILLCELL_X32 FILLCELL_168_1084 ();
 FILLCELL_X32 FILLCELL_168_1116 ();
 FILLCELL_X32 FILLCELL_168_1148 ();
 FILLCELL_X32 FILLCELL_168_1180 ();
 FILLCELL_X32 FILLCELL_168_1212 ();
 FILLCELL_X32 FILLCELL_168_1244 ();
 FILLCELL_X32 FILLCELL_168_1276 ();
 FILLCELL_X32 FILLCELL_168_1308 ();
 FILLCELL_X32 FILLCELL_168_1340 ();
 FILLCELL_X32 FILLCELL_168_1372 ();
 FILLCELL_X32 FILLCELL_168_1404 ();
 FILLCELL_X32 FILLCELL_168_1436 ();
 FILLCELL_X32 FILLCELL_168_1468 ();
 FILLCELL_X32 FILLCELL_168_1500 ();
 FILLCELL_X32 FILLCELL_168_1532 ();
 FILLCELL_X32 FILLCELL_168_1564 ();
 FILLCELL_X32 FILLCELL_168_1596 ();
 FILLCELL_X32 FILLCELL_168_1628 ();
 FILLCELL_X32 FILLCELL_168_1660 ();
 FILLCELL_X32 FILLCELL_168_1692 ();
 FILLCELL_X32 FILLCELL_168_1724 ();
 FILLCELL_X32 FILLCELL_168_1756 ();
 FILLCELL_X32 FILLCELL_168_1788 ();
 FILLCELL_X32 FILLCELL_168_1820 ();
 FILLCELL_X32 FILLCELL_168_1852 ();
 FILLCELL_X8 FILLCELL_168_1884 ();
 FILLCELL_X4 FILLCELL_168_1892 ();
 FILLCELL_X1 FILLCELL_168_1896 ();
 FILLCELL_X32 FILLCELL_169_0 ();
 FILLCELL_X32 FILLCELL_169_32 ();
 FILLCELL_X32 FILLCELL_169_64 ();
 FILLCELL_X32 FILLCELL_169_96 ();
 FILLCELL_X32 FILLCELL_169_128 ();
 FILLCELL_X16 FILLCELL_169_160 ();
 FILLCELL_X8 FILLCELL_169_176 ();
 FILLCELL_X4 FILLCELL_169_184 ();
 FILLCELL_X1 FILLCELL_169_188 ();
 FILLCELL_X32 FILLCELL_169_194 ();
 FILLCELL_X32 FILLCELL_169_226 ();
 FILLCELL_X32 FILLCELL_169_258 ();
 FILLCELL_X32 FILLCELL_169_290 ();
 FILLCELL_X32 FILLCELL_169_322 ();
 FILLCELL_X16 FILLCELL_169_354 ();
 FILLCELL_X8 FILLCELL_169_370 ();
 FILLCELL_X2 FILLCELL_169_378 ();
 FILLCELL_X1 FILLCELL_169_380 ();
 FILLCELL_X32 FILLCELL_169_384 ();
 FILLCELL_X32 FILLCELL_169_416 ();
 FILLCELL_X32 FILLCELL_169_448 ();
 FILLCELL_X32 FILLCELL_169_480 ();
 FILLCELL_X32 FILLCELL_169_512 ();
 FILLCELL_X32 FILLCELL_169_544 ();
 FILLCELL_X32 FILLCELL_169_576 ();
 FILLCELL_X32 FILLCELL_169_608 ();
 FILLCELL_X32 FILLCELL_169_640 ();
 FILLCELL_X32 FILLCELL_169_672 ();
 FILLCELL_X32 FILLCELL_169_704 ();
 FILLCELL_X32 FILLCELL_169_736 ();
 FILLCELL_X32 FILLCELL_169_768 ();
 FILLCELL_X32 FILLCELL_169_800 ();
 FILLCELL_X32 FILLCELL_169_832 ();
 FILLCELL_X32 FILLCELL_169_864 ();
 FILLCELL_X32 FILLCELL_169_896 ();
 FILLCELL_X32 FILLCELL_169_928 ();
 FILLCELL_X32 FILLCELL_169_960 ();
 FILLCELL_X32 FILLCELL_169_992 ();
 FILLCELL_X32 FILLCELL_169_1024 ();
 FILLCELL_X32 FILLCELL_169_1056 ();
 FILLCELL_X32 FILLCELL_169_1088 ();
 FILLCELL_X32 FILLCELL_169_1120 ();
 FILLCELL_X32 FILLCELL_169_1152 ();
 FILLCELL_X32 FILLCELL_169_1184 ();
 FILLCELL_X32 FILLCELL_169_1216 ();
 FILLCELL_X32 FILLCELL_169_1248 ();
 FILLCELL_X32 FILLCELL_169_1280 ();
 FILLCELL_X32 FILLCELL_169_1312 ();
 FILLCELL_X32 FILLCELL_169_1344 ();
 FILLCELL_X32 FILLCELL_169_1376 ();
 FILLCELL_X32 FILLCELL_169_1408 ();
 FILLCELL_X32 FILLCELL_169_1440 ();
 FILLCELL_X32 FILLCELL_169_1472 ();
 FILLCELL_X32 FILLCELL_169_1504 ();
 FILLCELL_X32 FILLCELL_169_1536 ();
 FILLCELL_X32 FILLCELL_169_1568 ();
 FILLCELL_X32 FILLCELL_169_1600 ();
 FILLCELL_X32 FILLCELL_169_1632 ();
 FILLCELL_X32 FILLCELL_169_1664 ();
 FILLCELL_X32 FILLCELL_169_1696 ();
 FILLCELL_X32 FILLCELL_169_1728 ();
 FILLCELL_X32 FILLCELL_169_1760 ();
 FILLCELL_X32 FILLCELL_169_1792 ();
 FILLCELL_X32 FILLCELL_169_1824 ();
 FILLCELL_X32 FILLCELL_169_1856 ();
 FILLCELL_X8 FILLCELL_169_1888 ();
 FILLCELL_X1 FILLCELL_169_1896 ();
 FILLCELL_X32 FILLCELL_170_0 ();
 FILLCELL_X32 FILLCELL_170_32 ();
 FILLCELL_X32 FILLCELL_170_64 ();
 FILLCELL_X32 FILLCELL_170_96 ();
 FILLCELL_X32 FILLCELL_170_128 ();
 FILLCELL_X16 FILLCELL_170_160 ();
 FILLCELL_X8 FILLCELL_170_176 ();
 FILLCELL_X32 FILLCELL_170_191 ();
 FILLCELL_X32 FILLCELL_170_223 ();
 FILLCELL_X32 FILLCELL_170_255 ();
 FILLCELL_X32 FILLCELL_170_287 ();
 FILLCELL_X32 FILLCELL_170_319 ();
 FILLCELL_X32 FILLCELL_170_351 ();
 FILLCELL_X32 FILLCELL_170_383 ();
 FILLCELL_X32 FILLCELL_170_415 ();
 FILLCELL_X32 FILLCELL_170_447 ();
 FILLCELL_X32 FILLCELL_170_479 ();
 FILLCELL_X32 FILLCELL_170_511 ();
 FILLCELL_X32 FILLCELL_170_543 ();
 FILLCELL_X32 FILLCELL_170_575 ();
 FILLCELL_X32 FILLCELL_170_607 ();
 FILLCELL_X32 FILLCELL_170_639 ();
 FILLCELL_X32 FILLCELL_170_671 ();
 FILLCELL_X32 FILLCELL_170_703 ();
 FILLCELL_X32 FILLCELL_170_735 ();
 FILLCELL_X32 FILLCELL_170_767 ();
 FILLCELL_X32 FILLCELL_170_799 ();
 FILLCELL_X32 FILLCELL_170_831 ();
 FILLCELL_X16 FILLCELL_170_863 ();
 FILLCELL_X8 FILLCELL_170_879 ();
 FILLCELL_X4 FILLCELL_170_887 ();
 FILLCELL_X2 FILLCELL_170_891 ();
 FILLCELL_X1 FILLCELL_170_893 ();
 FILLCELL_X32 FILLCELL_170_898 ();
 FILLCELL_X32 FILLCELL_170_930 ();
 FILLCELL_X32 FILLCELL_170_962 ();
 FILLCELL_X32 FILLCELL_170_994 ();
 FILLCELL_X32 FILLCELL_170_1026 ();
 FILLCELL_X32 FILLCELL_170_1058 ();
 FILLCELL_X32 FILLCELL_170_1090 ();
 FILLCELL_X32 FILLCELL_170_1122 ();
 FILLCELL_X32 FILLCELL_170_1154 ();
 FILLCELL_X32 FILLCELL_170_1186 ();
 FILLCELL_X32 FILLCELL_170_1218 ();
 FILLCELL_X32 FILLCELL_170_1250 ();
 FILLCELL_X32 FILLCELL_170_1282 ();
 FILLCELL_X32 FILLCELL_170_1314 ();
 FILLCELL_X32 FILLCELL_170_1346 ();
 FILLCELL_X32 FILLCELL_170_1378 ();
 FILLCELL_X32 FILLCELL_170_1410 ();
 FILLCELL_X32 FILLCELL_170_1442 ();
 FILLCELL_X32 FILLCELL_170_1474 ();
 FILLCELL_X32 FILLCELL_170_1506 ();
 FILLCELL_X32 FILLCELL_170_1538 ();
 FILLCELL_X32 FILLCELL_170_1570 ();
 FILLCELL_X32 FILLCELL_170_1602 ();
 FILLCELL_X32 FILLCELL_170_1634 ();
 FILLCELL_X32 FILLCELL_170_1666 ();
 FILLCELL_X32 FILLCELL_170_1698 ();
 FILLCELL_X32 FILLCELL_170_1730 ();
 FILLCELL_X32 FILLCELL_170_1762 ();
 FILLCELL_X32 FILLCELL_170_1794 ();
 FILLCELL_X32 FILLCELL_170_1826 ();
 FILLCELL_X32 FILLCELL_170_1858 ();
 FILLCELL_X4 FILLCELL_170_1890 ();
 FILLCELL_X2 FILLCELL_170_1894 ();
 FILLCELL_X1 FILLCELL_170_1896 ();
 FILLCELL_X32 FILLCELL_171_0 ();
 FILLCELL_X32 FILLCELL_171_32 ();
 FILLCELL_X32 FILLCELL_171_64 ();
 FILLCELL_X32 FILLCELL_171_96 ();
 FILLCELL_X32 FILLCELL_171_128 ();
 FILLCELL_X32 FILLCELL_171_160 ();
 FILLCELL_X32 FILLCELL_171_192 ();
 FILLCELL_X32 FILLCELL_171_224 ();
 FILLCELL_X32 FILLCELL_171_256 ();
 FILLCELL_X32 FILLCELL_171_288 ();
 FILLCELL_X32 FILLCELL_171_320 ();
 FILLCELL_X32 FILLCELL_171_352 ();
 FILLCELL_X32 FILLCELL_171_384 ();
 FILLCELL_X32 FILLCELL_171_416 ();
 FILLCELL_X32 FILLCELL_171_448 ();
 FILLCELL_X32 FILLCELL_171_480 ();
 FILLCELL_X32 FILLCELL_171_512 ();
 FILLCELL_X32 FILLCELL_171_544 ();
 FILLCELL_X32 FILLCELL_171_576 ();
 FILLCELL_X32 FILLCELL_171_608 ();
 FILLCELL_X32 FILLCELL_171_640 ();
 FILLCELL_X8 FILLCELL_171_672 ();
 FILLCELL_X2 FILLCELL_171_680 ();
 FILLCELL_X1 FILLCELL_171_682 ();
 FILLCELL_X32 FILLCELL_171_692 ();
 FILLCELL_X32 FILLCELL_171_724 ();
 FILLCELL_X32 FILLCELL_171_756 ();
 FILLCELL_X32 FILLCELL_171_788 ();
 FILLCELL_X32 FILLCELL_171_820 ();
 FILLCELL_X32 FILLCELL_171_852 ();
 FILLCELL_X32 FILLCELL_171_884 ();
 FILLCELL_X32 FILLCELL_171_916 ();
 FILLCELL_X32 FILLCELL_171_948 ();
 FILLCELL_X32 FILLCELL_171_980 ();
 FILLCELL_X32 FILLCELL_171_1012 ();
 FILLCELL_X32 FILLCELL_171_1044 ();
 FILLCELL_X32 FILLCELL_171_1076 ();
 FILLCELL_X32 FILLCELL_171_1108 ();
 FILLCELL_X32 FILLCELL_171_1140 ();
 FILLCELL_X32 FILLCELL_171_1172 ();
 FILLCELL_X32 FILLCELL_171_1204 ();
 FILLCELL_X32 FILLCELL_171_1236 ();
 FILLCELL_X32 FILLCELL_171_1268 ();
 FILLCELL_X32 FILLCELL_171_1300 ();
 FILLCELL_X32 FILLCELL_171_1332 ();
 FILLCELL_X32 FILLCELL_171_1364 ();
 FILLCELL_X32 FILLCELL_171_1396 ();
 FILLCELL_X32 FILLCELL_171_1428 ();
 FILLCELL_X32 FILLCELL_171_1460 ();
 FILLCELL_X32 FILLCELL_171_1492 ();
 FILLCELL_X32 FILLCELL_171_1524 ();
 FILLCELL_X32 FILLCELL_171_1556 ();
 FILLCELL_X32 FILLCELL_171_1588 ();
 FILLCELL_X32 FILLCELL_171_1620 ();
 FILLCELL_X32 FILLCELL_171_1652 ();
 FILLCELL_X32 FILLCELL_171_1684 ();
 FILLCELL_X32 FILLCELL_171_1716 ();
 FILLCELL_X32 FILLCELL_171_1748 ();
 FILLCELL_X32 FILLCELL_171_1780 ();
 FILLCELL_X32 FILLCELL_171_1812 ();
 FILLCELL_X32 FILLCELL_171_1844 ();
 FILLCELL_X16 FILLCELL_171_1876 ();
 FILLCELL_X4 FILLCELL_171_1892 ();
 FILLCELL_X1 FILLCELL_171_1896 ();
 FILLCELL_X32 FILLCELL_172_0 ();
 FILLCELL_X32 FILLCELL_172_32 ();
 FILLCELL_X32 FILLCELL_172_64 ();
 FILLCELL_X32 FILLCELL_172_96 ();
 FILLCELL_X32 FILLCELL_172_128 ();
 FILLCELL_X32 FILLCELL_172_160 ();
 FILLCELL_X32 FILLCELL_172_192 ();
 FILLCELL_X32 FILLCELL_172_224 ();
 FILLCELL_X32 FILLCELL_172_256 ();
 FILLCELL_X32 FILLCELL_172_288 ();
 FILLCELL_X32 FILLCELL_172_320 ();
 FILLCELL_X32 FILLCELL_172_352 ();
 FILLCELL_X32 FILLCELL_172_384 ();
 FILLCELL_X32 FILLCELL_172_416 ();
 FILLCELL_X32 FILLCELL_172_448 ();
 FILLCELL_X32 FILLCELL_172_480 ();
 FILLCELL_X32 FILLCELL_172_512 ();
 FILLCELL_X32 FILLCELL_172_544 ();
 FILLCELL_X32 FILLCELL_172_576 ();
 FILLCELL_X32 FILLCELL_172_608 ();
 FILLCELL_X32 FILLCELL_172_640 ();
 FILLCELL_X32 FILLCELL_172_672 ();
 FILLCELL_X32 FILLCELL_172_704 ();
 FILLCELL_X32 FILLCELL_172_736 ();
 FILLCELL_X32 FILLCELL_172_768 ();
 FILLCELL_X32 FILLCELL_172_800 ();
 FILLCELL_X32 FILLCELL_172_832 ();
 FILLCELL_X32 FILLCELL_172_864 ();
 FILLCELL_X32 FILLCELL_172_896 ();
 FILLCELL_X32 FILLCELL_172_928 ();
 FILLCELL_X32 FILLCELL_172_960 ();
 FILLCELL_X32 FILLCELL_172_992 ();
 FILLCELL_X32 FILLCELL_172_1024 ();
 FILLCELL_X32 FILLCELL_172_1056 ();
 FILLCELL_X32 FILLCELL_172_1088 ();
 FILLCELL_X32 FILLCELL_172_1120 ();
 FILLCELL_X32 FILLCELL_172_1152 ();
 FILLCELL_X32 FILLCELL_172_1184 ();
 FILLCELL_X32 FILLCELL_172_1216 ();
 FILLCELL_X32 FILLCELL_172_1248 ();
 FILLCELL_X32 FILLCELL_172_1280 ();
 FILLCELL_X32 FILLCELL_172_1312 ();
 FILLCELL_X32 FILLCELL_172_1344 ();
 FILLCELL_X32 FILLCELL_172_1376 ();
 FILLCELL_X32 FILLCELL_172_1408 ();
 FILLCELL_X32 FILLCELL_172_1440 ();
 FILLCELL_X32 FILLCELL_172_1472 ();
 FILLCELL_X32 FILLCELL_172_1504 ();
 FILLCELL_X32 FILLCELL_172_1536 ();
 FILLCELL_X32 FILLCELL_172_1568 ();
 FILLCELL_X32 FILLCELL_172_1600 ();
 FILLCELL_X32 FILLCELL_172_1632 ();
 FILLCELL_X32 FILLCELL_172_1664 ();
 FILLCELL_X32 FILLCELL_172_1696 ();
 FILLCELL_X32 FILLCELL_172_1728 ();
 FILLCELL_X32 FILLCELL_172_1760 ();
 FILLCELL_X32 FILLCELL_172_1792 ();
 FILLCELL_X32 FILLCELL_172_1824 ();
 FILLCELL_X32 FILLCELL_172_1856 ();
 FILLCELL_X8 FILLCELL_172_1888 ();
 FILLCELL_X1 FILLCELL_172_1896 ();
 FILLCELL_X32 FILLCELL_173_0 ();
 FILLCELL_X32 FILLCELL_173_32 ();
 FILLCELL_X32 FILLCELL_173_64 ();
 FILLCELL_X32 FILLCELL_173_96 ();
 FILLCELL_X32 FILLCELL_173_128 ();
 FILLCELL_X32 FILLCELL_173_160 ();
 FILLCELL_X32 FILLCELL_173_192 ();
 FILLCELL_X32 FILLCELL_173_224 ();
 FILLCELL_X32 FILLCELL_173_256 ();
 FILLCELL_X32 FILLCELL_173_292 ();
 FILLCELL_X32 FILLCELL_173_324 ();
 FILLCELL_X32 FILLCELL_173_356 ();
 FILLCELL_X32 FILLCELL_173_388 ();
 FILLCELL_X32 FILLCELL_173_420 ();
 FILLCELL_X32 FILLCELL_173_452 ();
 FILLCELL_X32 FILLCELL_173_484 ();
 FILLCELL_X32 FILLCELL_173_516 ();
 FILLCELL_X32 FILLCELL_173_548 ();
 FILLCELL_X32 FILLCELL_173_580 ();
 FILLCELL_X32 FILLCELL_173_612 ();
 FILLCELL_X32 FILLCELL_173_644 ();
 FILLCELL_X32 FILLCELL_173_676 ();
 FILLCELL_X32 FILLCELL_173_708 ();
 FILLCELL_X32 FILLCELL_173_740 ();
 FILLCELL_X32 FILLCELL_173_772 ();
 FILLCELL_X32 FILLCELL_173_804 ();
 FILLCELL_X32 FILLCELL_173_836 ();
 FILLCELL_X32 FILLCELL_173_868 ();
 FILLCELL_X8 FILLCELL_173_900 ();
 FILLCELL_X2 FILLCELL_173_908 ();
 FILLCELL_X32 FILLCELL_173_914 ();
 FILLCELL_X32 FILLCELL_173_946 ();
 FILLCELL_X32 FILLCELL_173_978 ();
 FILLCELL_X32 FILLCELL_173_1010 ();
 FILLCELL_X16 FILLCELL_173_1042 ();
 FILLCELL_X4 FILLCELL_173_1058 ();
 FILLCELL_X32 FILLCELL_173_1066 ();
 FILLCELL_X32 FILLCELL_173_1098 ();
 FILLCELL_X32 FILLCELL_173_1130 ();
 FILLCELL_X32 FILLCELL_173_1162 ();
 FILLCELL_X32 FILLCELL_173_1194 ();
 FILLCELL_X32 FILLCELL_173_1226 ();
 FILLCELL_X32 FILLCELL_173_1258 ();
 FILLCELL_X32 FILLCELL_173_1290 ();
 FILLCELL_X32 FILLCELL_173_1322 ();
 FILLCELL_X32 FILLCELL_173_1354 ();
 FILLCELL_X32 FILLCELL_173_1386 ();
 FILLCELL_X32 FILLCELL_173_1418 ();
 FILLCELL_X32 FILLCELL_173_1450 ();
 FILLCELL_X32 FILLCELL_173_1482 ();
 FILLCELL_X32 FILLCELL_173_1514 ();
 FILLCELL_X32 FILLCELL_173_1546 ();
 FILLCELL_X32 FILLCELL_173_1578 ();
 FILLCELL_X32 FILLCELL_173_1610 ();
 FILLCELL_X32 FILLCELL_173_1642 ();
 FILLCELL_X32 FILLCELL_173_1674 ();
 FILLCELL_X32 FILLCELL_173_1706 ();
 FILLCELL_X32 FILLCELL_173_1738 ();
 FILLCELL_X32 FILLCELL_173_1770 ();
 FILLCELL_X32 FILLCELL_173_1802 ();
 FILLCELL_X32 FILLCELL_173_1834 ();
 FILLCELL_X16 FILLCELL_173_1866 ();
 FILLCELL_X8 FILLCELL_173_1882 ();
 FILLCELL_X4 FILLCELL_173_1890 ();
 FILLCELL_X2 FILLCELL_173_1894 ();
 FILLCELL_X1 FILLCELL_173_1896 ();
 FILLCELL_X32 FILLCELL_174_0 ();
 FILLCELL_X32 FILLCELL_174_32 ();
 FILLCELL_X32 FILLCELL_174_64 ();
 FILLCELL_X32 FILLCELL_174_96 ();
 FILLCELL_X32 FILLCELL_174_128 ();
 FILLCELL_X32 FILLCELL_174_160 ();
 FILLCELL_X32 FILLCELL_174_192 ();
 FILLCELL_X32 FILLCELL_174_224 ();
 FILLCELL_X32 FILLCELL_174_256 ();
 FILLCELL_X32 FILLCELL_174_288 ();
 FILLCELL_X16 FILLCELL_174_320 ();
 FILLCELL_X8 FILLCELL_174_336 ();
 FILLCELL_X4 FILLCELL_174_344 ();
 FILLCELL_X2 FILLCELL_174_348 ();
 FILLCELL_X1 FILLCELL_174_350 ();
 FILLCELL_X32 FILLCELL_174_355 ();
 FILLCELL_X32 FILLCELL_174_387 ();
 FILLCELL_X32 FILLCELL_174_419 ();
 FILLCELL_X32 FILLCELL_174_451 ();
 FILLCELL_X32 FILLCELL_174_483 ();
 FILLCELL_X32 FILLCELL_174_515 ();
 FILLCELL_X16 FILLCELL_174_547 ();
 FILLCELL_X2 FILLCELL_174_563 ();
 FILLCELL_X1 FILLCELL_174_565 ();
 FILLCELL_X32 FILLCELL_174_575 ();
 FILLCELL_X32 FILLCELL_174_607 ();
 FILLCELL_X8 FILLCELL_174_639 ();
 FILLCELL_X1 FILLCELL_174_647 ();
 FILLCELL_X32 FILLCELL_174_654 ();
 FILLCELL_X32 FILLCELL_174_686 ();
 FILLCELL_X32 FILLCELL_174_718 ();
 FILLCELL_X1 FILLCELL_174_750 ();
 FILLCELL_X32 FILLCELL_174_755 ();
 FILLCELL_X32 FILLCELL_174_787 ();
 FILLCELL_X32 FILLCELL_174_819 ();
 FILLCELL_X32 FILLCELL_174_851 ();
 FILLCELL_X32 FILLCELL_174_883 ();
 FILLCELL_X32 FILLCELL_174_915 ();
 FILLCELL_X32 FILLCELL_174_947 ();
 FILLCELL_X32 FILLCELL_174_979 ();
 FILLCELL_X2 FILLCELL_174_1011 ();
 FILLCELL_X32 FILLCELL_174_1016 ();
 FILLCELL_X32 FILLCELL_174_1048 ();
 FILLCELL_X32 FILLCELL_174_1080 ();
 FILLCELL_X32 FILLCELL_174_1112 ();
 FILLCELL_X32 FILLCELL_174_1144 ();
 FILLCELL_X32 FILLCELL_174_1176 ();
 FILLCELL_X32 FILLCELL_174_1208 ();
 FILLCELL_X32 FILLCELL_174_1240 ();
 FILLCELL_X32 FILLCELL_174_1272 ();
 FILLCELL_X32 FILLCELL_174_1304 ();
 FILLCELL_X32 FILLCELL_174_1336 ();
 FILLCELL_X32 FILLCELL_174_1368 ();
 FILLCELL_X32 FILLCELL_174_1400 ();
 FILLCELL_X32 FILLCELL_174_1432 ();
 FILLCELL_X32 FILLCELL_174_1464 ();
 FILLCELL_X32 FILLCELL_174_1496 ();
 FILLCELL_X32 FILLCELL_174_1528 ();
 FILLCELL_X32 FILLCELL_174_1560 ();
 FILLCELL_X32 FILLCELL_174_1592 ();
 FILLCELL_X32 FILLCELL_174_1624 ();
 FILLCELL_X32 FILLCELL_174_1656 ();
 FILLCELL_X32 FILLCELL_174_1688 ();
 FILLCELL_X32 FILLCELL_174_1720 ();
 FILLCELL_X32 FILLCELL_174_1752 ();
 FILLCELL_X32 FILLCELL_174_1784 ();
 FILLCELL_X32 FILLCELL_174_1816 ();
 FILLCELL_X32 FILLCELL_174_1848 ();
 FILLCELL_X16 FILLCELL_174_1880 ();
 FILLCELL_X1 FILLCELL_174_1896 ();
 FILLCELL_X32 FILLCELL_175_0 ();
 FILLCELL_X32 FILLCELL_175_32 ();
 FILLCELL_X32 FILLCELL_175_64 ();
 FILLCELL_X32 FILLCELL_175_96 ();
 FILLCELL_X32 FILLCELL_175_128 ();
 FILLCELL_X32 FILLCELL_175_160 ();
 FILLCELL_X32 FILLCELL_175_192 ();
 FILLCELL_X32 FILLCELL_175_224 ();
 FILLCELL_X32 FILLCELL_175_256 ();
 FILLCELL_X32 FILLCELL_175_288 ();
 FILLCELL_X32 FILLCELL_175_320 ();
 FILLCELL_X32 FILLCELL_175_352 ();
 FILLCELL_X32 FILLCELL_175_384 ();
 FILLCELL_X32 FILLCELL_175_416 ();
 FILLCELL_X32 FILLCELL_175_448 ();
 FILLCELL_X32 FILLCELL_175_480 ();
 FILLCELL_X32 FILLCELL_175_512 ();
 FILLCELL_X32 FILLCELL_175_544 ();
 FILLCELL_X32 FILLCELL_175_576 ();
 FILLCELL_X32 FILLCELL_175_608 ();
 FILLCELL_X32 FILLCELL_175_640 ();
 FILLCELL_X32 FILLCELL_175_672 ();
 FILLCELL_X32 FILLCELL_175_704 ();
 FILLCELL_X16 FILLCELL_175_736 ();
 FILLCELL_X8 FILLCELL_175_752 ();
 FILLCELL_X4 FILLCELL_175_760 ();
 FILLCELL_X2 FILLCELL_175_764 ();
 FILLCELL_X1 FILLCELL_175_766 ();
 FILLCELL_X32 FILLCELL_175_772 ();
 FILLCELL_X32 FILLCELL_175_804 ();
 FILLCELL_X32 FILLCELL_175_836 ();
 FILLCELL_X32 FILLCELL_175_868 ();
 FILLCELL_X32 FILLCELL_175_900 ();
 FILLCELL_X32 FILLCELL_175_932 ();
 FILLCELL_X8 FILLCELL_175_964 ();
 FILLCELL_X32 FILLCELL_175_977 ();
 FILLCELL_X32 FILLCELL_175_1012 ();
 FILLCELL_X32 FILLCELL_175_1044 ();
 FILLCELL_X32 FILLCELL_175_1076 ();
 FILLCELL_X32 FILLCELL_175_1108 ();
 FILLCELL_X32 FILLCELL_175_1140 ();
 FILLCELL_X32 FILLCELL_175_1172 ();
 FILLCELL_X32 FILLCELL_175_1204 ();
 FILLCELL_X32 FILLCELL_175_1236 ();
 FILLCELL_X32 FILLCELL_175_1268 ();
 FILLCELL_X32 FILLCELL_175_1300 ();
 FILLCELL_X32 FILLCELL_175_1332 ();
 FILLCELL_X32 FILLCELL_175_1364 ();
 FILLCELL_X32 FILLCELL_175_1396 ();
 FILLCELL_X32 FILLCELL_175_1428 ();
 FILLCELL_X32 FILLCELL_175_1460 ();
 FILLCELL_X32 FILLCELL_175_1492 ();
 FILLCELL_X32 FILLCELL_175_1524 ();
 FILLCELL_X32 FILLCELL_175_1556 ();
 FILLCELL_X32 FILLCELL_175_1588 ();
 FILLCELL_X32 FILLCELL_175_1620 ();
 FILLCELL_X32 FILLCELL_175_1652 ();
 FILLCELL_X32 FILLCELL_175_1684 ();
 FILLCELL_X32 FILLCELL_175_1716 ();
 FILLCELL_X32 FILLCELL_175_1748 ();
 FILLCELL_X32 FILLCELL_175_1780 ();
 FILLCELL_X32 FILLCELL_175_1812 ();
 FILLCELL_X32 FILLCELL_175_1844 ();
 FILLCELL_X16 FILLCELL_175_1876 ();
 FILLCELL_X4 FILLCELL_175_1892 ();
 FILLCELL_X1 FILLCELL_175_1896 ();
 FILLCELL_X32 FILLCELL_176_0 ();
 FILLCELL_X32 FILLCELL_176_32 ();
 FILLCELL_X32 FILLCELL_176_64 ();
 FILLCELL_X32 FILLCELL_176_96 ();
 FILLCELL_X32 FILLCELL_176_128 ();
 FILLCELL_X32 FILLCELL_176_160 ();
 FILLCELL_X32 FILLCELL_176_192 ();
 FILLCELL_X32 FILLCELL_176_224 ();
 FILLCELL_X32 FILLCELL_176_256 ();
 FILLCELL_X32 FILLCELL_176_288 ();
 FILLCELL_X32 FILLCELL_176_320 ();
 FILLCELL_X32 FILLCELL_176_352 ();
 FILLCELL_X32 FILLCELL_176_384 ();
 FILLCELL_X32 FILLCELL_176_416 ();
 FILLCELL_X32 FILLCELL_176_448 ();
 FILLCELL_X32 FILLCELL_176_480 ();
 FILLCELL_X32 FILLCELL_176_512 ();
 FILLCELL_X32 FILLCELL_176_544 ();
 FILLCELL_X32 FILLCELL_176_576 ();
 FILLCELL_X32 FILLCELL_176_608 ();
 FILLCELL_X32 FILLCELL_176_640 ();
 FILLCELL_X32 FILLCELL_176_672 ();
 FILLCELL_X32 FILLCELL_176_704 ();
 FILLCELL_X32 FILLCELL_176_736 ();
 FILLCELL_X32 FILLCELL_176_768 ();
 FILLCELL_X32 FILLCELL_176_800 ();
 FILLCELL_X32 FILLCELL_176_832 ();
 FILLCELL_X32 FILLCELL_176_864 ();
 FILLCELL_X32 FILLCELL_176_896 ();
 FILLCELL_X32 FILLCELL_176_928 ();
 FILLCELL_X32 FILLCELL_176_960 ();
 FILLCELL_X32 FILLCELL_176_992 ();
 FILLCELL_X32 FILLCELL_176_1024 ();
 FILLCELL_X8 FILLCELL_176_1056 ();
 FILLCELL_X4 FILLCELL_176_1064 ();
 FILLCELL_X2 FILLCELL_176_1068 ();
 FILLCELL_X32 FILLCELL_176_1075 ();
 FILLCELL_X32 FILLCELL_176_1107 ();
 FILLCELL_X32 FILLCELL_176_1139 ();
 FILLCELL_X32 FILLCELL_176_1171 ();
 FILLCELL_X32 FILLCELL_176_1203 ();
 FILLCELL_X32 FILLCELL_176_1235 ();
 FILLCELL_X32 FILLCELL_176_1267 ();
 FILLCELL_X32 FILLCELL_176_1299 ();
 FILLCELL_X32 FILLCELL_176_1331 ();
 FILLCELL_X32 FILLCELL_176_1363 ();
 FILLCELL_X32 FILLCELL_176_1395 ();
 FILLCELL_X32 FILLCELL_176_1427 ();
 FILLCELL_X32 FILLCELL_176_1459 ();
 FILLCELL_X32 FILLCELL_176_1491 ();
 FILLCELL_X32 FILLCELL_176_1523 ();
 FILLCELL_X32 FILLCELL_176_1555 ();
 FILLCELL_X32 FILLCELL_176_1587 ();
 FILLCELL_X32 FILLCELL_176_1619 ();
 FILLCELL_X32 FILLCELL_176_1651 ();
 FILLCELL_X32 FILLCELL_176_1683 ();
 FILLCELL_X32 FILLCELL_176_1715 ();
 FILLCELL_X32 FILLCELL_176_1747 ();
 FILLCELL_X32 FILLCELL_176_1779 ();
 FILLCELL_X32 FILLCELL_176_1811 ();
 FILLCELL_X32 FILLCELL_176_1843 ();
 FILLCELL_X16 FILLCELL_176_1875 ();
 FILLCELL_X4 FILLCELL_176_1891 ();
 FILLCELL_X2 FILLCELL_176_1895 ();
 FILLCELL_X32 FILLCELL_177_0 ();
 FILLCELL_X32 FILLCELL_177_32 ();
 FILLCELL_X32 FILLCELL_177_64 ();
 FILLCELL_X32 FILLCELL_177_96 ();
 FILLCELL_X32 FILLCELL_177_128 ();
 FILLCELL_X32 FILLCELL_177_160 ();
 FILLCELL_X32 FILLCELL_177_192 ();
 FILLCELL_X32 FILLCELL_177_224 ();
 FILLCELL_X16 FILLCELL_177_256 ();
 FILLCELL_X8 FILLCELL_177_272 ();
 FILLCELL_X2 FILLCELL_177_280 ();
 FILLCELL_X32 FILLCELL_177_286 ();
 FILLCELL_X32 FILLCELL_177_318 ();
 FILLCELL_X8 FILLCELL_177_350 ();
 FILLCELL_X4 FILLCELL_177_358 ();
 FILLCELL_X32 FILLCELL_177_366 ();
 FILLCELL_X32 FILLCELL_177_398 ();
 FILLCELL_X32 FILLCELL_177_430 ();
 FILLCELL_X32 FILLCELL_177_462 ();
 FILLCELL_X32 FILLCELL_177_494 ();
 FILLCELL_X32 FILLCELL_177_526 ();
 FILLCELL_X32 FILLCELL_177_558 ();
 FILLCELL_X32 FILLCELL_177_590 ();
 FILLCELL_X32 FILLCELL_177_622 ();
 FILLCELL_X32 FILLCELL_177_654 ();
 FILLCELL_X32 FILLCELL_177_686 ();
 FILLCELL_X32 FILLCELL_177_718 ();
 FILLCELL_X16 FILLCELL_177_750 ();
 FILLCELL_X2 FILLCELL_177_766 ();
 FILLCELL_X32 FILLCELL_177_772 ();
 FILLCELL_X32 FILLCELL_177_804 ();
 FILLCELL_X32 FILLCELL_177_836 ();
 FILLCELL_X32 FILLCELL_177_868 ();
 FILLCELL_X16 FILLCELL_177_900 ();
 FILLCELL_X32 FILLCELL_177_920 ();
 FILLCELL_X16 FILLCELL_177_952 ();
 FILLCELL_X8 FILLCELL_177_968 ();
 FILLCELL_X2 FILLCELL_177_976 ();
 FILLCELL_X32 FILLCELL_177_981 ();
 FILLCELL_X16 FILLCELL_177_1013 ();
 FILLCELL_X8 FILLCELL_177_1029 ();
 FILLCELL_X4 FILLCELL_177_1037 ();
 FILLCELL_X32 FILLCELL_177_1043 ();
 FILLCELL_X32 FILLCELL_177_1075 ();
 FILLCELL_X32 FILLCELL_177_1107 ();
 FILLCELL_X32 FILLCELL_177_1139 ();
 FILLCELL_X32 FILLCELL_177_1171 ();
 FILLCELL_X32 FILLCELL_177_1203 ();
 FILLCELL_X32 FILLCELL_177_1235 ();
 FILLCELL_X32 FILLCELL_177_1267 ();
 FILLCELL_X32 FILLCELL_177_1299 ();
 FILLCELL_X32 FILLCELL_177_1331 ();
 FILLCELL_X32 FILLCELL_177_1363 ();
 FILLCELL_X32 FILLCELL_177_1395 ();
 FILLCELL_X32 FILLCELL_177_1427 ();
 FILLCELL_X32 FILLCELL_177_1459 ();
 FILLCELL_X32 FILLCELL_177_1491 ();
 FILLCELL_X32 FILLCELL_177_1523 ();
 FILLCELL_X32 FILLCELL_177_1555 ();
 FILLCELL_X32 FILLCELL_177_1587 ();
 FILLCELL_X32 FILLCELL_177_1619 ();
 FILLCELL_X32 FILLCELL_177_1651 ();
 FILLCELL_X32 FILLCELL_177_1683 ();
 FILLCELL_X32 FILLCELL_177_1715 ();
 FILLCELL_X32 FILLCELL_177_1747 ();
 FILLCELL_X32 FILLCELL_177_1779 ();
 FILLCELL_X32 FILLCELL_177_1811 ();
 FILLCELL_X32 FILLCELL_177_1843 ();
 FILLCELL_X16 FILLCELL_177_1875 ();
 FILLCELL_X4 FILLCELL_177_1891 ();
 FILLCELL_X2 FILLCELL_177_1895 ();
 FILLCELL_X32 FILLCELL_178_0 ();
 FILLCELL_X32 FILLCELL_178_32 ();
 FILLCELL_X32 FILLCELL_178_64 ();
 FILLCELL_X32 FILLCELL_178_96 ();
 FILLCELL_X32 FILLCELL_178_128 ();
 FILLCELL_X32 FILLCELL_178_160 ();
 FILLCELL_X32 FILLCELL_178_192 ();
 FILLCELL_X32 FILLCELL_178_224 ();
 FILLCELL_X32 FILLCELL_178_256 ();
 FILLCELL_X32 FILLCELL_178_288 ();
 FILLCELL_X32 FILLCELL_178_320 ();
 FILLCELL_X32 FILLCELL_178_352 ();
 FILLCELL_X32 FILLCELL_178_384 ();
 FILLCELL_X32 FILLCELL_178_416 ();
 FILLCELL_X4 FILLCELL_178_448 ();
 FILLCELL_X2 FILLCELL_178_452 ();
 FILLCELL_X32 FILLCELL_178_459 ();
 FILLCELL_X32 FILLCELL_178_491 ();
 FILLCELL_X32 FILLCELL_178_523 ();
 FILLCELL_X32 FILLCELL_178_555 ();
 FILLCELL_X32 FILLCELL_178_587 ();
 FILLCELL_X32 FILLCELL_178_619 ();
 FILLCELL_X32 FILLCELL_178_651 ();
 FILLCELL_X32 FILLCELL_178_683 ();
 FILLCELL_X32 FILLCELL_178_715 ();
 FILLCELL_X32 FILLCELL_178_747 ();
 FILLCELL_X32 FILLCELL_178_779 ();
 FILLCELL_X32 FILLCELL_178_811 ();
 FILLCELL_X32 FILLCELL_178_843 ();
 FILLCELL_X32 FILLCELL_178_875 ();
 FILLCELL_X32 FILLCELL_178_907 ();
 FILLCELL_X32 FILLCELL_178_939 ();
 FILLCELL_X16 FILLCELL_178_971 ();
 FILLCELL_X8 FILLCELL_178_987 ();
 FILLCELL_X4 FILLCELL_178_995 ();
 FILLCELL_X1 FILLCELL_178_999 ();
 FILLCELL_X32 FILLCELL_178_1002 ();
 FILLCELL_X32 FILLCELL_178_1034 ();
 FILLCELL_X8 FILLCELL_178_1066 ();
 FILLCELL_X4 FILLCELL_178_1074 ();
 FILLCELL_X1 FILLCELL_178_1078 ();
 FILLCELL_X32 FILLCELL_178_1086 ();
 FILLCELL_X32 FILLCELL_178_1118 ();
 FILLCELL_X32 FILLCELL_178_1150 ();
 FILLCELL_X32 FILLCELL_178_1182 ();
 FILLCELL_X32 FILLCELL_178_1214 ();
 FILLCELL_X32 FILLCELL_178_1246 ();
 FILLCELL_X32 FILLCELL_178_1278 ();
 FILLCELL_X32 FILLCELL_178_1310 ();
 FILLCELL_X32 FILLCELL_178_1342 ();
 FILLCELL_X32 FILLCELL_178_1374 ();
 FILLCELL_X32 FILLCELL_178_1406 ();
 FILLCELL_X32 FILLCELL_178_1438 ();
 FILLCELL_X32 FILLCELL_178_1470 ();
 FILLCELL_X32 FILLCELL_178_1502 ();
 FILLCELL_X32 FILLCELL_178_1534 ();
 FILLCELL_X32 FILLCELL_178_1566 ();
 FILLCELL_X32 FILLCELL_178_1598 ();
 FILLCELL_X32 FILLCELL_178_1630 ();
 FILLCELL_X32 FILLCELL_178_1662 ();
 FILLCELL_X32 FILLCELL_178_1694 ();
 FILLCELL_X32 FILLCELL_178_1726 ();
 FILLCELL_X32 FILLCELL_178_1758 ();
 FILLCELL_X32 FILLCELL_178_1790 ();
 FILLCELL_X32 FILLCELL_178_1822 ();
 FILLCELL_X32 FILLCELL_178_1854 ();
 FILLCELL_X8 FILLCELL_178_1886 ();
 FILLCELL_X2 FILLCELL_178_1894 ();
 FILLCELL_X1 FILLCELL_178_1896 ();
 FILLCELL_X32 FILLCELL_179_0 ();
 FILLCELL_X32 FILLCELL_179_32 ();
 FILLCELL_X32 FILLCELL_179_64 ();
 FILLCELL_X32 FILLCELL_179_96 ();
 FILLCELL_X32 FILLCELL_179_128 ();
 FILLCELL_X32 FILLCELL_179_160 ();
 FILLCELL_X32 FILLCELL_179_192 ();
 FILLCELL_X32 FILLCELL_179_224 ();
 FILLCELL_X32 FILLCELL_179_256 ();
 FILLCELL_X32 FILLCELL_179_288 ();
 FILLCELL_X32 FILLCELL_179_320 ();
 FILLCELL_X4 FILLCELL_179_352 ();
 FILLCELL_X2 FILLCELL_179_356 ();
 FILLCELL_X32 FILLCELL_179_361 ();
 FILLCELL_X32 FILLCELL_179_393 ();
 FILLCELL_X32 FILLCELL_179_425 ();
 FILLCELL_X32 FILLCELL_179_457 ();
 FILLCELL_X16 FILLCELL_179_489 ();
 FILLCELL_X8 FILLCELL_179_505 ();
 FILLCELL_X2 FILLCELL_179_513 ();
 FILLCELL_X1 FILLCELL_179_515 ();
 FILLCELL_X32 FILLCELL_179_519 ();
 FILLCELL_X32 FILLCELL_179_551 ();
 FILLCELL_X32 FILLCELL_179_583 ();
 FILLCELL_X32 FILLCELL_179_615 ();
 FILLCELL_X32 FILLCELL_179_647 ();
 FILLCELL_X32 FILLCELL_179_679 ();
 FILLCELL_X32 FILLCELL_179_711 ();
 FILLCELL_X32 FILLCELL_179_743 ();
 FILLCELL_X8 FILLCELL_179_775 ();
 FILLCELL_X4 FILLCELL_179_783 ();
 FILLCELL_X2 FILLCELL_179_787 ();
 FILLCELL_X1 FILLCELL_179_789 ();
 FILLCELL_X32 FILLCELL_179_793 ();
 FILLCELL_X32 FILLCELL_179_825 ();
 FILLCELL_X32 FILLCELL_179_857 ();
 FILLCELL_X32 FILLCELL_179_889 ();
 FILLCELL_X32 FILLCELL_179_921 ();
 FILLCELL_X32 FILLCELL_179_953 ();
 FILLCELL_X32 FILLCELL_179_985 ();
 FILLCELL_X32 FILLCELL_179_1017 ();
 FILLCELL_X32 FILLCELL_179_1049 ();
 FILLCELL_X32 FILLCELL_179_1081 ();
 FILLCELL_X32 FILLCELL_179_1113 ();
 FILLCELL_X32 FILLCELL_179_1145 ();
 FILLCELL_X32 FILLCELL_179_1177 ();
 FILLCELL_X32 FILLCELL_179_1209 ();
 FILLCELL_X32 FILLCELL_179_1241 ();
 FILLCELL_X32 FILLCELL_179_1273 ();
 FILLCELL_X32 FILLCELL_179_1305 ();
 FILLCELL_X32 FILLCELL_179_1337 ();
 FILLCELL_X32 FILLCELL_179_1369 ();
 FILLCELL_X32 FILLCELL_179_1401 ();
 FILLCELL_X32 FILLCELL_179_1433 ();
 FILLCELL_X32 FILLCELL_179_1465 ();
 FILLCELL_X32 FILLCELL_179_1497 ();
 FILLCELL_X32 FILLCELL_179_1529 ();
 FILLCELL_X32 FILLCELL_179_1561 ();
 FILLCELL_X32 FILLCELL_179_1593 ();
 FILLCELL_X32 FILLCELL_179_1625 ();
 FILLCELL_X32 FILLCELL_179_1657 ();
 FILLCELL_X32 FILLCELL_179_1689 ();
 FILLCELL_X32 FILLCELL_179_1721 ();
 FILLCELL_X32 FILLCELL_179_1753 ();
 FILLCELL_X32 FILLCELL_179_1785 ();
 FILLCELL_X32 FILLCELL_179_1817 ();
 FILLCELL_X32 FILLCELL_179_1849 ();
 FILLCELL_X16 FILLCELL_179_1881 ();
 FILLCELL_X32 FILLCELL_180_0 ();
 FILLCELL_X32 FILLCELL_180_32 ();
 FILLCELL_X32 FILLCELL_180_64 ();
 FILLCELL_X32 FILLCELL_180_96 ();
 FILLCELL_X32 FILLCELL_180_128 ();
 FILLCELL_X32 FILLCELL_180_160 ();
 FILLCELL_X32 FILLCELL_180_192 ();
 FILLCELL_X16 FILLCELL_180_224 ();
 FILLCELL_X8 FILLCELL_180_240 ();
 FILLCELL_X2 FILLCELL_180_248 ();
 FILLCELL_X32 FILLCELL_180_253 ();
 FILLCELL_X32 FILLCELL_180_285 ();
 FILLCELL_X32 FILLCELL_180_317 ();
 FILLCELL_X32 FILLCELL_180_349 ();
 FILLCELL_X32 FILLCELL_180_381 ();
 FILLCELL_X32 FILLCELL_180_413 ();
 FILLCELL_X32 FILLCELL_180_445 ();
 FILLCELL_X32 FILLCELL_180_477 ();
 FILLCELL_X32 FILLCELL_180_509 ();
 FILLCELL_X32 FILLCELL_180_541 ();
 FILLCELL_X32 FILLCELL_180_573 ();
 FILLCELL_X32 FILLCELL_180_605 ();
 FILLCELL_X32 FILLCELL_180_637 ();
 FILLCELL_X32 FILLCELL_180_669 ();
 FILLCELL_X32 FILLCELL_180_701 ();
 FILLCELL_X32 FILLCELL_180_733 ();
 FILLCELL_X32 FILLCELL_180_765 ();
 FILLCELL_X32 FILLCELL_180_797 ();
 FILLCELL_X32 FILLCELL_180_829 ();
 FILLCELL_X32 FILLCELL_180_861 ();
 FILLCELL_X32 FILLCELL_180_893 ();
 FILLCELL_X32 FILLCELL_180_925 ();
 FILLCELL_X32 FILLCELL_180_957 ();
 FILLCELL_X32 FILLCELL_180_989 ();
 FILLCELL_X32 FILLCELL_180_1021 ();
 FILLCELL_X32 FILLCELL_180_1053 ();
 FILLCELL_X32 FILLCELL_180_1085 ();
 FILLCELL_X4 FILLCELL_180_1117 ();
 FILLCELL_X32 FILLCELL_180_1138 ();
 FILLCELL_X32 FILLCELL_180_1170 ();
 FILLCELL_X32 FILLCELL_180_1202 ();
 FILLCELL_X32 FILLCELL_180_1234 ();
 FILLCELL_X32 FILLCELL_180_1266 ();
 FILLCELL_X32 FILLCELL_180_1298 ();
 FILLCELL_X32 FILLCELL_180_1330 ();
 FILLCELL_X32 FILLCELL_180_1362 ();
 FILLCELL_X32 FILLCELL_180_1394 ();
 FILLCELL_X32 FILLCELL_180_1426 ();
 FILLCELL_X32 FILLCELL_180_1458 ();
 FILLCELL_X32 FILLCELL_180_1490 ();
 FILLCELL_X32 FILLCELL_180_1522 ();
 FILLCELL_X32 FILLCELL_180_1554 ();
 FILLCELL_X32 FILLCELL_180_1586 ();
 FILLCELL_X32 FILLCELL_180_1618 ();
 FILLCELL_X32 FILLCELL_180_1650 ();
 FILLCELL_X32 FILLCELL_180_1682 ();
 FILLCELL_X32 FILLCELL_180_1714 ();
 FILLCELL_X32 FILLCELL_180_1746 ();
 FILLCELL_X32 FILLCELL_180_1778 ();
 FILLCELL_X32 FILLCELL_180_1810 ();
 FILLCELL_X32 FILLCELL_180_1842 ();
 FILLCELL_X16 FILLCELL_180_1874 ();
 FILLCELL_X4 FILLCELL_180_1890 ();
 FILLCELL_X2 FILLCELL_180_1894 ();
 FILLCELL_X1 FILLCELL_180_1896 ();
 FILLCELL_X32 FILLCELL_181_0 ();
 FILLCELL_X32 FILLCELL_181_32 ();
 FILLCELL_X32 FILLCELL_181_64 ();
 FILLCELL_X32 FILLCELL_181_96 ();
 FILLCELL_X32 FILLCELL_181_128 ();
 FILLCELL_X32 FILLCELL_181_160 ();
 FILLCELL_X32 FILLCELL_181_192 ();
 FILLCELL_X32 FILLCELL_181_224 ();
 FILLCELL_X32 FILLCELL_181_256 ();
 FILLCELL_X32 FILLCELL_181_288 ();
 FILLCELL_X32 FILLCELL_181_320 ();
 FILLCELL_X32 FILLCELL_181_352 ();
 FILLCELL_X32 FILLCELL_181_384 ();
 FILLCELL_X32 FILLCELL_181_416 ();
 FILLCELL_X32 FILLCELL_181_448 ();
 FILLCELL_X32 FILLCELL_181_480 ();
 FILLCELL_X8 FILLCELL_181_512 ();
 FILLCELL_X2 FILLCELL_181_520 ();
 FILLCELL_X1 FILLCELL_181_522 ();
 FILLCELL_X32 FILLCELL_181_526 ();
 FILLCELL_X4 FILLCELL_181_558 ();
 FILLCELL_X2 FILLCELL_181_562 ();
 FILLCELL_X1 FILLCELL_181_564 ();
 FILLCELL_X32 FILLCELL_181_570 ();
 FILLCELL_X32 FILLCELL_181_602 ();
 FILLCELL_X32 FILLCELL_181_634 ();
 FILLCELL_X32 FILLCELL_181_666 ();
 FILLCELL_X32 FILLCELL_181_698 ();
 FILLCELL_X32 FILLCELL_181_730 ();
 FILLCELL_X32 FILLCELL_181_762 ();
 FILLCELL_X32 FILLCELL_181_794 ();
 FILLCELL_X32 FILLCELL_181_826 ();
 FILLCELL_X16 FILLCELL_181_858 ();
 FILLCELL_X32 FILLCELL_181_878 ();
 FILLCELL_X8 FILLCELL_181_910 ();
 FILLCELL_X4 FILLCELL_181_918 ();
 FILLCELL_X1 FILLCELL_181_922 ();
 FILLCELL_X32 FILLCELL_181_926 ();
 FILLCELL_X32 FILLCELL_181_958 ();
 FILLCELL_X32 FILLCELL_181_990 ();
 FILLCELL_X32 FILLCELL_181_1022 ();
 FILLCELL_X32 FILLCELL_181_1054 ();
 FILLCELL_X32 FILLCELL_181_1086 ();
 FILLCELL_X32 FILLCELL_181_1118 ();
 FILLCELL_X32 FILLCELL_181_1150 ();
 FILLCELL_X32 FILLCELL_181_1182 ();
 FILLCELL_X32 FILLCELL_181_1214 ();
 FILLCELL_X32 FILLCELL_181_1246 ();
 FILLCELL_X32 FILLCELL_181_1278 ();
 FILLCELL_X32 FILLCELL_181_1310 ();
 FILLCELL_X32 FILLCELL_181_1342 ();
 FILLCELL_X32 FILLCELL_181_1374 ();
 FILLCELL_X32 FILLCELL_181_1406 ();
 FILLCELL_X32 FILLCELL_181_1438 ();
 FILLCELL_X32 FILLCELL_181_1470 ();
 FILLCELL_X32 FILLCELL_181_1502 ();
 FILLCELL_X32 FILLCELL_181_1534 ();
 FILLCELL_X32 FILLCELL_181_1566 ();
 FILLCELL_X32 FILLCELL_181_1598 ();
 FILLCELL_X32 FILLCELL_181_1630 ();
 FILLCELL_X32 FILLCELL_181_1662 ();
 FILLCELL_X32 FILLCELL_181_1694 ();
 FILLCELL_X32 FILLCELL_181_1726 ();
 FILLCELL_X32 FILLCELL_181_1758 ();
 FILLCELL_X32 FILLCELL_181_1790 ();
 FILLCELL_X32 FILLCELL_181_1822 ();
 FILLCELL_X32 FILLCELL_181_1854 ();
 FILLCELL_X8 FILLCELL_181_1886 ();
 FILLCELL_X2 FILLCELL_181_1894 ();
 FILLCELL_X1 FILLCELL_181_1896 ();
 FILLCELL_X32 FILLCELL_182_0 ();
 FILLCELL_X32 FILLCELL_182_32 ();
 FILLCELL_X32 FILLCELL_182_64 ();
 FILLCELL_X32 FILLCELL_182_96 ();
 FILLCELL_X32 FILLCELL_182_128 ();
 FILLCELL_X32 FILLCELL_182_160 ();
 FILLCELL_X32 FILLCELL_182_192 ();
 FILLCELL_X32 FILLCELL_182_224 ();
 FILLCELL_X32 FILLCELL_182_256 ();
 FILLCELL_X32 FILLCELL_182_288 ();
 FILLCELL_X32 FILLCELL_182_320 ();
 FILLCELL_X8 FILLCELL_182_352 ();
 FILLCELL_X2 FILLCELL_182_360 ();
 FILLCELL_X1 FILLCELL_182_362 ();
 FILLCELL_X32 FILLCELL_182_366 ();
 FILLCELL_X32 FILLCELL_182_398 ();
 FILLCELL_X8 FILLCELL_182_430 ();
 FILLCELL_X4 FILLCELL_182_438 ();
 FILLCELL_X1 FILLCELL_182_442 ();
 FILLCELL_X32 FILLCELL_182_447 ();
 FILLCELL_X32 FILLCELL_182_479 ();
 FILLCELL_X32 FILLCELL_182_511 ();
 FILLCELL_X8 FILLCELL_182_543 ();
 FILLCELL_X4 FILLCELL_182_551 ();
 FILLCELL_X2 FILLCELL_182_555 ();
 FILLCELL_X1 FILLCELL_182_557 ();
 FILLCELL_X32 FILLCELL_182_563 ();
 FILLCELL_X32 FILLCELL_182_595 ();
 FILLCELL_X32 FILLCELL_182_627 ();
 FILLCELL_X16 FILLCELL_182_659 ();
 FILLCELL_X4 FILLCELL_182_675 ();
 FILLCELL_X1 FILLCELL_182_679 ();
 FILLCELL_X16 FILLCELL_182_683 ();
 FILLCELL_X1 FILLCELL_182_699 ();
 FILLCELL_X32 FILLCELL_182_703 ();
 FILLCELL_X32 FILLCELL_182_735 ();
 FILLCELL_X32 FILLCELL_182_767 ();
 FILLCELL_X16 FILLCELL_182_799 ();
 FILLCELL_X8 FILLCELL_182_815 ();
 FILLCELL_X4 FILLCELL_182_823 ();
 FILLCELL_X32 FILLCELL_182_830 ();
 FILLCELL_X32 FILLCELL_182_862 ();
 FILLCELL_X32 FILLCELL_182_894 ();
 FILLCELL_X32 FILLCELL_182_926 ();
 FILLCELL_X32 FILLCELL_182_958 ();
 FILLCELL_X32 FILLCELL_182_990 ();
 FILLCELL_X32 FILLCELL_182_1022 ();
 FILLCELL_X32 FILLCELL_182_1054 ();
 FILLCELL_X32 FILLCELL_182_1086 ();
 FILLCELL_X32 FILLCELL_182_1118 ();
 FILLCELL_X32 FILLCELL_182_1150 ();
 FILLCELL_X32 FILLCELL_182_1182 ();
 FILLCELL_X32 FILLCELL_182_1214 ();
 FILLCELL_X32 FILLCELL_182_1246 ();
 FILLCELL_X32 FILLCELL_182_1278 ();
 FILLCELL_X32 FILLCELL_182_1310 ();
 FILLCELL_X32 FILLCELL_182_1342 ();
 FILLCELL_X32 FILLCELL_182_1374 ();
 FILLCELL_X32 FILLCELL_182_1406 ();
 FILLCELL_X32 FILLCELL_182_1438 ();
 FILLCELL_X32 FILLCELL_182_1470 ();
 FILLCELL_X32 FILLCELL_182_1502 ();
 FILLCELL_X32 FILLCELL_182_1534 ();
 FILLCELL_X32 FILLCELL_182_1566 ();
 FILLCELL_X32 FILLCELL_182_1598 ();
 FILLCELL_X32 FILLCELL_182_1630 ();
 FILLCELL_X32 FILLCELL_182_1662 ();
 FILLCELL_X32 FILLCELL_182_1694 ();
 FILLCELL_X32 FILLCELL_182_1726 ();
 FILLCELL_X32 FILLCELL_182_1758 ();
 FILLCELL_X32 FILLCELL_182_1790 ();
 FILLCELL_X32 FILLCELL_182_1822 ();
 FILLCELL_X32 FILLCELL_182_1854 ();
 FILLCELL_X8 FILLCELL_182_1886 ();
 FILLCELL_X2 FILLCELL_182_1894 ();
 FILLCELL_X1 FILLCELL_182_1896 ();
 FILLCELL_X32 FILLCELL_183_0 ();
 FILLCELL_X32 FILLCELL_183_32 ();
 FILLCELL_X32 FILLCELL_183_64 ();
 FILLCELL_X32 FILLCELL_183_96 ();
 FILLCELL_X32 FILLCELL_183_128 ();
 FILLCELL_X32 FILLCELL_183_160 ();
 FILLCELL_X32 FILLCELL_183_192 ();
 FILLCELL_X32 FILLCELL_183_224 ();
 FILLCELL_X32 FILLCELL_183_256 ();
 FILLCELL_X32 FILLCELL_183_288 ();
 FILLCELL_X32 FILLCELL_183_320 ();
 FILLCELL_X32 FILLCELL_183_352 ();
 FILLCELL_X32 FILLCELL_183_384 ();
 FILLCELL_X32 FILLCELL_183_416 ();
 FILLCELL_X2 FILLCELL_183_448 ();
 FILLCELL_X32 FILLCELL_183_455 ();
 FILLCELL_X32 FILLCELL_183_487 ();
 FILLCELL_X32 FILLCELL_183_519 ();
 FILLCELL_X16 FILLCELL_183_551 ();
 FILLCELL_X8 FILLCELL_183_567 ();
 FILLCELL_X32 FILLCELL_183_578 ();
 FILLCELL_X32 FILLCELL_183_610 ();
 FILLCELL_X32 FILLCELL_183_642 ();
 FILLCELL_X32 FILLCELL_183_674 ();
 FILLCELL_X32 FILLCELL_183_706 ();
 FILLCELL_X32 FILLCELL_183_738 ();
 FILLCELL_X32 FILLCELL_183_770 ();
 FILLCELL_X32 FILLCELL_183_802 ();
 FILLCELL_X32 FILLCELL_183_834 ();
 FILLCELL_X32 FILLCELL_183_866 ();
 FILLCELL_X32 FILLCELL_183_898 ();
 FILLCELL_X32 FILLCELL_183_930 ();
 FILLCELL_X32 FILLCELL_183_962 ();
 FILLCELL_X32 FILLCELL_183_994 ();
 FILLCELL_X32 FILLCELL_183_1026 ();
 FILLCELL_X32 FILLCELL_183_1058 ();
 FILLCELL_X32 FILLCELL_183_1090 ();
 FILLCELL_X32 FILLCELL_183_1122 ();
 FILLCELL_X32 FILLCELL_183_1154 ();
 FILLCELL_X32 FILLCELL_183_1186 ();
 FILLCELL_X32 FILLCELL_183_1218 ();
 FILLCELL_X32 FILLCELL_183_1250 ();
 FILLCELL_X32 FILLCELL_183_1282 ();
 FILLCELL_X32 FILLCELL_183_1314 ();
 FILLCELL_X32 FILLCELL_183_1346 ();
 FILLCELL_X32 FILLCELL_183_1378 ();
 FILLCELL_X32 FILLCELL_183_1410 ();
 FILLCELL_X32 FILLCELL_183_1442 ();
 FILLCELL_X32 FILLCELL_183_1474 ();
 FILLCELL_X32 FILLCELL_183_1506 ();
 FILLCELL_X32 FILLCELL_183_1538 ();
 FILLCELL_X32 FILLCELL_183_1570 ();
 FILLCELL_X32 FILLCELL_183_1602 ();
 FILLCELL_X32 FILLCELL_183_1634 ();
 FILLCELL_X32 FILLCELL_183_1666 ();
 FILLCELL_X32 FILLCELL_183_1698 ();
 FILLCELL_X32 FILLCELL_183_1730 ();
 FILLCELL_X32 FILLCELL_183_1762 ();
 FILLCELL_X32 FILLCELL_183_1794 ();
 FILLCELL_X32 FILLCELL_183_1826 ();
 FILLCELL_X32 FILLCELL_183_1858 ();
 FILLCELL_X4 FILLCELL_183_1890 ();
 FILLCELL_X2 FILLCELL_183_1894 ();
 FILLCELL_X1 FILLCELL_183_1896 ();
 FILLCELL_X32 FILLCELL_184_0 ();
 FILLCELL_X32 FILLCELL_184_32 ();
 FILLCELL_X32 FILLCELL_184_64 ();
 FILLCELL_X32 FILLCELL_184_96 ();
 FILLCELL_X16 FILLCELL_184_128 ();
 FILLCELL_X8 FILLCELL_184_144 ();
 FILLCELL_X4 FILLCELL_184_152 ();
 FILLCELL_X1 FILLCELL_184_156 ();
 FILLCELL_X32 FILLCELL_184_160 ();
 FILLCELL_X32 FILLCELL_184_192 ();
 FILLCELL_X32 FILLCELL_184_224 ();
 FILLCELL_X32 FILLCELL_184_256 ();
 FILLCELL_X32 FILLCELL_184_288 ();
 FILLCELL_X32 FILLCELL_184_320 ();
 FILLCELL_X32 FILLCELL_184_352 ();
 FILLCELL_X32 FILLCELL_184_384 ();
 FILLCELL_X16 FILLCELL_184_416 ();
 FILLCELL_X8 FILLCELL_184_432 ();
 FILLCELL_X32 FILLCELL_184_444 ();
 FILLCELL_X32 FILLCELL_184_476 ();
 FILLCELL_X32 FILLCELL_184_508 ();
 FILLCELL_X32 FILLCELL_184_540 ();
 FILLCELL_X32 FILLCELL_184_572 ();
 FILLCELL_X32 FILLCELL_184_604 ();
 FILLCELL_X32 FILLCELL_184_636 ();
 FILLCELL_X2 FILLCELL_184_668 ();
 FILLCELL_X32 FILLCELL_184_679 ();
 FILLCELL_X32 FILLCELL_184_711 ();
 FILLCELL_X32 FILLCELL_184_743 ();
 FILLCELL_X32 FILLCELL_184_775 ();
 FILLCELL_X32 FILLCELL_184_807 ();
 FILLCELL_X16 FILLCELL_184_839 ();
 FILLCELL_X8 FILLCELL_184_855 ();
 FILLCELL_X32 FILLCELL_184_867 ();
 FILLCELL_X32 FILLCELL_184_899 ();
 FILLCELL_X32 FILLCELL_184_931 ();
 FILLCELL_X32 FILLCELL_184_963 ();
 FILLCELL_X32 FILLCELL_184_995 ();
 FILLCELL_X32 FILLCELL_184_1027 ();
 FILLCELL_X32 FILLCELL_184_1059 ();
 FILLCELL_X32 FILLCELL_184_1091 ();
 FILLCELL_X32 FILLCELL_184_1123 ();
 FILLCELL_X32 FILLCELL_184_1155 ();
 FILLCELL_X32 FILLCELL_184_1187 ();
 FILLCELL_X32 FILLCELL_184_1219 ();
 FILLCELL_X32 FILLCELL_184_1251 ();
 FILLCELL_X32 FILLCELL_184_1283 ();
 FILLCELL_X32 FILLCELL_184_1315 ();
 FILLCELL_X32 FILLCELL_184_1347 ();
 FILLCELL_X32 FILLCELL_184_1379 ();
 FILLCELL_X32 FILLCELL_184_1411 ();
 FILLCELL_X32 FILLCELL_184_1443 ();
 FILLCELL_X32 FILLCELL_184_1475 ();
 FILLCELL_X32 FILLCELL_184_1507 ();
 FILLCELL_X32 FILLCELL_184_1539 ();
 FILLCELL_X32 FILLCELL_184_1571 ();
 FILLCELL_X32 FILLCELL_184_1603 ();
 FILLCELL_X32 FILLCELL_184_1635 ();
 FILLCELL_X32 FILLCELL_184_1667 ();
 FILLCELL_X32 FILLCELL_184_1699 ();
 FILLCELL_X32 FILLCELL_184_1731 ();
 FILLCELL_X32 FILLCELL_184_1763 ();
 FILLCELL_X32 FILLCELL_184_1795 ();
 FILLCELL_X32 FILLCELL_184_1827 ();
 FILLCELL_X32 FILLCELL_184_1859 ();
 FILLCELL_X4 FILLCELL_184_1891 ();
 FILLCELL_X2 FILLCELL_184_1895 ();
 FILLCELL_X32 FILLCELL_185_0 ();
 FILLCELL_X32 FILLCELL_185_32 ();
 FILLCELL_X32 FILLCELL_185_64 ();
 FILLCELL_X32 FILLCELL_185_96 ();
 FILLCELL_X32 FILLCELL_185_128 ();
 FILLCELL_X32 FILLCELL_185_160 ();
 FILLCELL_X32 FILLCELL_185_192 ();
 FILLCELL_X8 FILLCELL_185_224 ();
 FILLCELL_X32 FILLCELL_185_235 ();
 FILLCELL_X32 FILLCELL_185_267 ();
 FILLCELL_X32 FILLCELL_185_299 ();
 FILLCELL_X32 FILLCELL_185_331 ();
 FILLCELL_X32 FILLCELL_185_363 ();
 FILLCELL_X32 FILLCELL_185_395 ();
 FILLCELL_X32 FILLCELL_185_427 ();
 FILLCELL_X32 FILLCELL_185_459 ();
 FILLCELL_X32 FILLCELL_185_491 ();
 FILLCELL_X32 FILLCELL_185_523 ();
 FILLCELL_X32 FILLCELL_185_555 ();
 FILLCELL_X32 FILLCELL_185_587 ();
 FILLCELL_X32 FILLCELL_185_619 ();
 FILLCELL_X32 FILLCELL_185_651 ();
 FILLCELL_X32 FILLCELL_185_683 ();
 FILLCELL_X16 FILLCELL_185_715 ();
 FILLCELL_X8 FILLCELL_185_731 ();
 FILLCELL_X4 FILLCELL_185_739 ();
 FILLCELL_X1 FILLCELL_185_743 ();
 FILLCELL_X32 FILLCELL_185_749 ();
 FILLCELL_X32 FILLCELL_185_781 ();
 FILLCELL_X32 FILLCELL_185_813 ();
 FILLCELL_X32 FILLCELL_185_845 ();
 FILLCELL_X32 FILLCELL_185_877 ();
 FILLCELL_X32 FILLCELL_185_909 ();
 FILLCELL_X32 FILLCELL_185_941 ();
 FILLCELL_X32 FILLCELL_185_973 ();
 FILLCELL_X32 FILLCELL_185_1005 ();
 FILLCELL_X32 FILLCELL_185_1037 ();
 FILLCELL_X32 FILLCELL_185_1069 ();
 FILLCELL_X32 FILLCELL_185_1101 ();
 FILLCELL_X32 FILLCELL_185_1133 ();
 FILLCELL_X32 FILLCELL_185_1165 ();
 FILLCELL_X32 FILLCELL_185_1197 ();
 FILLCELL_X32 FILLCELL_185_1229 ();
 FILLCELL_X32 FILLCELL_185_1261 ();
 FILLCELL_X32 FILLCELL_185_1293 ();
 FILLCELL_X32 FILLCELL_185_1325 ();
 FILLCELL_X32 FILLCELL_185_1357 ();
 FILLCELL_X32 FILLCELL_185_1389 ();
 FILLCELL_X32 FILLCELL_185_1421 ();
 FILLCELL_X32 FILLCELL_185_1453 ();
 FILLCELL_X32 FILLCELL_185_1485 ();
 FILLCELL_X32 FILLCELL_185_1517 ();
 FILLCELL_X32 FILLCELL_185_1549 ();
 FILLCELL_X32 FILLCELL_185_1581 ();
 FILLCELL_X32 FILLCELL_185_1613 ();
 FILLCELL_X32 FILLCELL_185_1645 ();
 FILLCELL_X32 FILLCELL_185_1677 ();
 FILLCELL_X32 FILLCELL_185_1709 ();
 FILLCELL_X32 FILLCELL_185_1741 ();
 FILLCELL_X32 FILLCELL_185_1773 ();
 FILLCELL_X32 FILLCELL_185_1805 ();
 FILLCELL_X32 FILLCELL_185_1837 ();
 FILLCELL_X16 FILLCELL_185_1869 ();
 FILLCELL_X8 FILLCELL_185_1885 ();
 FILLCELL_X4 FILLCELL_185_1893 ();
 FILLCELL_X32 FILLCELL_186_0 ();
 FILLCELL_X32 FILLCELL_186_32 ();
 FILLCELL_X32 FILLCELL_186_64 ();
 FILLCELL_X32 FILLCELL_186_96 ();
 FILLCELL_X32 FILLCELL_186_128 ();
 FILLCELL_X32 FILLCELL_186_160 ();
 FILLCELL_X16 FILLCELL_186_192 ();
 FILLCELL_X8 FILLCELL_186_208 ();
 FILLCELL_X2 FILLCELL_186_216 ();
 FILLCELL_X1 FILLCELL_186_218 ();
 FILLCELL_X32 FILLCELL_186_236 ();
 FILLCELL_X32 FILLCELL_186_268 ();
 FILLCELL_X32 FILLCELL_186_300 ();
 FILLCELL_X32 FILLCELL_186_332 ();
 FILLCELL_X32 FILLCELL_186_364 ();
 FILLCELL_X32 FILLCELL_186_396 ();
 FILLCELL_X32 FILLCELL_186_428 ();
 FILLCELL_X32 FILLCELL_186_460 ();
 FILLCELL_X32 FILLCELL_186_492 ();
 FILLCELL_X8 FILLCELL_186_524 ();
 FILLCELL_X32 FILLCELL_186_537 ();
 FILLCELL_X32 FILLCELL_186_569 ();
 FILLCELL_X32 FILLCELL_186_601 ();
 FILLCELL_X32 FILLCELL_186_633 ();
 FILLCELL_X32 FILLCELL_186_665 ();
 FILLCELL_X32 FILLCELL_186_697 ();
 FILLCELL_X32 FILLCELL_186_729 ();
 FILLCELL_X32 FILLCELL_186_761 ();
 FILLCELL_X16 FILLCELL_186_793 ();
 FILLCELL_X8 FILLCELL_186_809 ();
 FILLCELL_X4 FILLCELL_186_817 ();
 FILLCELL_X2 FILLCELL_186_821 ();
 FILLCELL_X1 FILLCELL_186_823 ();
 FILLCELL_X32 FILLCELL_186_841 ();
 FILLCELL_X32 FILLCELL_186_873 ();
 FILLCELL_X32 FILLCELL_186_905 ();
 FILLCELL_X32 FILLCELL_186_937 ();
 FILLCELL_X32 FILLCELL_186_969 ();
 FILLCELL_X32 FILLCELL_186_1001 ();
 FILLCELL_X32 FILLCELL_186_1033 ();
 FILLCELL_X32 FILLCELL_186_1065 ();
 FILLCELL_X32 FILLCELL_186_1097 ();
 FILLCELL_X32 FILLCELL_186_1129 ();
 FILLCELL_X32 FILLCELL_186_1161 ();
 FILLCELL_X32 FILLCELL_186_1193 ();
 FILLCELL_X32 FILLCELL_186_1225 ();
 FILLCELL_X32 FILLCELL_186_1257 ();
 FILLCELL_X32 FILLCELL_186_1289 ();
 FILLCELL_X32 FILLCELL_186_1321 ();
 FILLCELL_X32 FILLCELL_186_1353 ();
 FILLCELL_X32 FILLCELL_186_1385 ();
 FILLCELL_X32 FILLCELL_186_1417 ();
 FILLCELL_X32 FILLCELL_186_1449 ();
 FILLCELL_X32 FILLCELL_186_1481 ();
 FILLCELL_X32 FILLCELL_186_1513 ();
 FILLCELL_X32 FILLCELL_186_1545 ();
 FILLCELL_X32 FILLCELL_186_1577 ();
 FILLCELL_X32 FILLCELL_186_1609 ();
 FILLCELL_X32 FILLCELL_186_1641 ();
 FILLCELL_X32 FILLCELL_186_1673 ();
 FILLCELL_X32 FILLCELL_186_1705 ();
 FILLCELL_X32 FILLCELL_186_1737 ();
 FILLCELL_X32 FILLCELL_186_1769 ();
 FILLCELL_X32 FILLCELL_186_1801 ();
 FILLCELL_X32 FILLCELL_186_1833 ();
 FILLCELL_X32 FILLCELL_186_1865 ();
 FILLCELL_X32 FILLCELL_187_0 ();
 FILLCELL_X32 FILLCELL_187_32 ();
 FILLCELL_X32 FILLCELL_187_64 ();
 FILLCELL_X32 FILLCELL_187_96 ();
 FILLCELL_X32 FILLCELL_187_128 ();
 FILLCELL_X32 FILLCELL_187_160 ();
 FILLCELL_X32 FILLCELL_187_192 ();
 FILLCELL_X32 FILLCELL_187_224 ();
 FILLCELL_X4 FILLCELL_187_256 ();
 FILLCELL_X32 FILLCELL_187_264 ();
 FILLCELL_X32 FILLCELL_187_296 ();
 FILLCELL_X16 FILLCELL_187_328 ();
 FILLCELL_X1 FILLCELL_187_344 ();
 FILLCELL_X32 FILLCELL_187_362 ();
 FILLCELL_X32 FILLCELL_187_394 ();
 FILLCELL_X32 FILLCELL_187_426 ();
 FILLCELL_X32 FILLCELL_187_458 ();
 FILLCELL_X32 FILLCELL_187_490 ();
 FILLCELL_X32 FILLCELL_187_522 ();
 FILLCELL_X32 FILLCELL_187_554 ();
 FILLCELL_X32 FILLCELL_187_586 ();
 FILLCELL_X32 FILLCELL_187_618 ();
 FILLCELL_X32 FILLCELL_187_650 ();
 FILLCELL_X32 FILLCELL_187_682 ();
 FILLCELL_X32 FILLCELL_187_714 ();
 FILLCELL_X32 FILLCELL_187_746 ();
 FILLCELL_X32 FILLCELL_187_778 ();
 FILLCELL_X32 FILLCELL_187_810 ();
 FILLCELL_X32 FILLCELL_187_842 ();
 FILLCELL_X32 FILLCELL_187_874 ();
 FILLCELL_X32 FILLCELL_187_906 ();
 FILLCELL_X32 FILLCELL_187_938 ();
 FILLCELL_X32 FILLCELL_187_970 ();
 FILLCELL_X32 FILLCELL_187_1002 ();
 FILLCELL_X32 FILLCELL_187_1034 ();
 FILLCELL_X32 FILLCELL_187_1066 ();
 FILLCELL_X32 FILLCELL_187_1098 ();
 FILLCELL_X32 FILLCELL_187_1130 ();
 FILLCELL_X32 FILLCELL_187_1162 ();
 FILLCELL_X32 FILLCELL_187_1194 ();
 FILLCELL_X32 FILLCELL_187_1226 ();
 FILLCELL_X32 FILLCELL_187_1258 ();
 FILLCELL_X32 FILLCELL_187_1290 ();
 FILLCELL_X32 FILLCELL_187_1322 ();
 FILLCELL_X32 FILLCELL_187_1354 ();
 FILLCELL_X32 FILLCELL_187_1386 ();
 FILLCELL_X32 FILLCELL_187_1418 ();
 FILLCELL_X32 FILLCELL_187_1450 ();
 FILLCELL_X32 FILLCELL_187_1482 ();
 FILLCELL_X32 FILLCELL_187_1514 ();
 FILLCELL_X32 FILLCELL_187_1546 ();
 FILLCELL_X32 FILLCELL_187_1578 ();
 FILLCELL_X32 FILLCELL_187_1610 ();
 FILLCELL_X32 FILLCELL_187_1642 ();
 FILLCELL_X32 FILLCELL_187_1674 ();
 FILLCELL_X32 FILLCELL_187_1706 ();
 FILLCELL_X32 FILLCELL_187_1738 ();
 FILLCELL_X32 FILLCELL_187_1770 ();
 FILLCELL_X32 FILLCELL_187_1802 ();
 FILLCELL_X32 FILLCELL_187_1834 ();
 FILLCELL_X16 FILLCELL_187_1866 ();
 FILLCELL_X8 FILLCELL_187_1882 ();
 FILLCELL_X4 FILLCELL_187_1890 ();
 FILLCELL_X2 FILLCELL_187_1894 ();
 FILLCELL_X1 FILLCELL_187_1896 ();
 FILLCELL_X32 FILLCELL_188_0 ();
 FILLCELL_X32 FILLCELL_188_32 ();
 FILLCELL_X32 FILLCELL_188_64 ();
 FILLCELL_X32 FILLCELL_188_96 ();
 FILLCELL_X32 FILLCELL_188_128 ();
 FILLCELL_X32 FILLCELL_188_160 ();
 FILLCELL_X32 FILLCELL_188_192 ();
 FILLCELL_X4 FILLCELL_188_224 ();
 FILLCELL_X32 FILLCELL_188_232 ();
 FILLCELL_X32 FILLCELL_188_264 ();
 FILLCELL_X32 FILLCELL_188_296 ();
 FILLCELL_X32 FILLCELL_188_328 ();
 FILLCELL_X32 FILLCELL_188_360 ();
 FILLCELL_X32 FILLCELL_188_392 ();
 FILLCELL_X32 FILLCELL_188_424 ();
 FILLCELL_X32 FILLCELL_188_456 ();
 FILLCELL_X32 FILLCELL_188_488 ();
 FILLCELL_X32 FILLCELL_188_520 ();
 FILLCELL_X32 FILLCELL_188_552 ();
 FILLCELL_X32 FILLCELL_188_584 ();
 FILLCELL_X32 FILLCELL_188_616 ();
 FILLCELL_X32 FILLCELL_188_648 ();
 FILLCELL_X32 FILLCELL_188_680 ();
 FILLCELL_X32 FILLCELL_188_712 ();
 FILLCELL_X32 FILLCELL_188_744 ();
 FILLCELL_X32 FILLCELL_188_776 ();
 FILLCELL_X32 FILLCELL_188_808 ();
 FILLCELL_X32 FILLCELL_188_840 ();
 FILLCELL_X32 FILLCELL_188_872 ();
 FILLCELL_X32 FILLCELL_188_904 ();
 FILLCELL_X8 FILLCELL_188_936 ();
 FILLCELL_X4 FILLCELL_188_944 ();
 FILLCELL_X2 FILLCELL_188_948 ();
 FILLCELL_X1 FILLCELL_188_950 ();
 FILLCELL_X32 FILLCELL_188_955 ();
 FILLCELL_X32 FILLCELL_188_987 ();
 FILLCELL_X32 FILLCELL_188_1019 ();
 FILLCELL_X32 FILLCELL_188_1051 ();
 FILLCELL_X32 FILLCELL_188_1083 ();
 FILLCELL_X32 FILLCELL_188_1115 ();
 FILLCELL_X32 FILLCELL_188_1147 ();
 FILLCELL_X32 FILLCELL_188_1179 ();
 FILLCELL_X32 FILLCELL_188_1211 ();
 FILLCELL_X32 FILLCELL_188_1243 ();
 FILLCELL_X32 FILLCELL_188_1275 ();
 FILLCELL_X32 FILLCELL_188_1307 ();
 FILLCELL_X32 FILLCELL_188_1339 ();
 FILLCELL_X32 FILLCELL_188_1371 ();
 FILLCELL_X32 FILLCELL_188_1403 ();
 FILLCELL_X32 FILLCELL_188_1435 ();
 FILLCELL_X32 FILLCELL_188_1467 ();
 FILLCELL_X32 FILLCELL_188_1499 ();
 FILLCELL_X32 FILLCELL_188_1531 ();
 FILLCELL_X32 FILLCELL_188_1563 ();
 FILLCELL_X32 FILLCELL_188_1595 ();
 FILLCELL_X32 FILLCELL_188_1627 ();
 FILLCELL_X32 FILLCELL_188_1659 ();
 FILLCELL_X32 FILLCELL_188_1691 ();
 FILLCELL_X32 FILLCELL_188_1723 ();
 FILLCELL_X32 FILLCELL_188_1755 ();
 FILLCELL_X32 FILLCELL_188_1787 ();
 FILLCELL_X32 FILLCELL_188_1819 ();
 FILLCELL_X32 FILLCELL_188_1851 ();
 FILLCELL_X8 FILLCELL_188_1883 ();
 FILLCELL_X4 FILLCELL_188_1891 ();
 FILLCELL_X2 FILLCELL_188_1895 ();
 FILLCELL_X32 FILLCELL_189_0 ();
 FILLCELL_X32 FILLCELL_189_32 ();
 FILLCELL_X32 FILLCELL_189_64 ();
 FILLCELL_X32 FILLCELL_189_96 ();
 FILLCELL_X32 FILLCELL_189_128 ();
 FILLCELL_X32 FILLCELL_189_160 ();
 FILLCELL_X32 FILLCELL_189_192 ();
 FILLCELL_X32 FILLCELL_189_224 ();
 FILLCELL_X32 FILLCELL_189_256 ();
 FILLCELL_X32 FILLCELL_189_288 ();
 FILLCELL_X32 FILLCELL_189_320 ();
 FILLCELL_X32 FILLCELL_189_352 ();
 FILLCELL_X32 FILLCELL_189_384 ();
 FILLCELL_X32 FILLCELL_189_416 ();
 FILLCELL_X32 FILLCELL_189_448 ();
 FILLCELL_X32 FILLCELL_189_480 ();
 FILLCELL_X32 FILLCELL_189_512 ();
 FILLCELL_X32 FILLCELL_189_544 ();
 FILLCELL_X32 FILLCELL_189_576 ();
 FILLCELL_X32 FILLCELL_189_608 ();
 FILLCELL_X32 FILLCELL_189_640 ();
 FILLCELL_X32 FILLCELL_189_672 ();
 FILLCELL_X32 FILLCELL_189_704 ();
 FILLCELL_X32 FILLCELL_189_736 ();
 FILLCELL_X32 FILLCELL_189_768 ();
 FILLCELL_X32 FILLCELL_189_800 ();
 FILLCELL_X32 FILLCELL_189_832 ();
 FILLCELL_X32 FILLCELL_189_864 ();
 FILLCELL_X16 FILLCELL_189_896 ();
 FILLCELL_X8 FILLCELL_189_912 ();
 FILLCELL_X4 FILLCELL_189_920 ();
 FILLCELL_X2 FILLCELL_189_924 ();
 FILLCELL_X1 FILLCELL_189_926 ();
 FILLCELL_X8 FILLCELL_189_931 ();
 FILLCELL_X2 FILLCELL_189_939 ();
 FILLCELL_X32 FILLCELL_189_944 ();
 FILLCELL_X32 FILLCELL_189_976 ();
 FILLCELL_X32 FILLCELL_189_1008 ();
 FILLCELL_X32 FILLCELL_189_1040 ();
 FILLCELL_X32 FILLCELL_189_1072 ();
 FILLCELL_X32 FILLCELL_189_1104 ();
 FILLCELL_X32 FILLCELL_189_1136 ();
 FILLCELL_X32 FILLCELL_189_1168 ();
 FILLCELL_X32 FILLCELL_189_1200 ();
 FILLCELL_X32 FILLCELL_189_1232 ();
 FILLCELL_X32 FILLCELL_189_1264 ();
 FILLCELL_X32 FILLCELL_189_1296 ();
 FILLCELL_X32 FILLCELL_189_1328 ();
 FILLCELL_X32 FILLCELL_189_1360 ();
 FILLCELL_X32 FILLCELL_189_1392 ();
 FILLCELL_X32 FILLCELL_189_1424 ();
 FILLCELL_X32 FILLCELL_189_1456 ();
 FILLCELL_X32 FILLCELL_189_1488 ();
 FILLCELL_X32 FILLCELL_189_1520 ();
 FILLCELL_X32 FILLCELL_189_1552 ();
 FILLCELL_X32 FILLCELL_189_1584 ();
 FILLCELL_X32 FILLCELL_189_1616 ();
 FILLCELL_X32 FILLCELL_189_1648 ();
 FILLCELL_X32 FILLCELL_189_1680 ();
 FILLCELL_X32 FILLCELL_189_1712 ();
 FILLCELL_X32 FILLCELL_189_1744 ();
 FILLCELL_X32 FILLCELL_189_1776 ();
 FILLCELL_X32 FILLCELL_189_1808 ();
 FILLCELL_X32 FILLCELL_189_1840 ();
 FILLCELL_X16 FILLCELL_189_1872 ();
 FILLCELL_X8 FILLCELL_189_1888 ();
 FILLCELL_X1 FILLCELL_189_1896 ();
 FILLCELL_X32 FILLCELL_190_0 ();
 FILLCELL_X32 FILLCELL_190_32 ();
 FILLCELL_X32 FILLCELL_190_64 ();
 FILLCELL_X32 FILLCELL_190_96 ();
 FILLCELL_X32 FILLCELL_190_128 ();
 FILLCELL_X32 FILLCELL_190_160 ();
 FILLCELL_X32 FILLCELL_190_192 ();
 FILLCELL_X32 FILLCELL_190_224 ();
 FILLCELL_X32 FILLCELL_190_256 ();
 FILLCELL_X32 FILLCELL_190_288 ();
 FILLCELL_X32 FILLCELL_190_320 ();
 FILLCELL_X32 FILLCELL_190_352 ();
 FILLCELL_X8 FILLCELL_190_384 ();
 FILLCELL_X4 FILLCELL_190_392 ();
 FILLCELL_X32 FILLCELL_190_398 ();
 FILLCELL_X32 FILLCELL_190_430 ();
 FILLCELL_X32 FILLCELL_190_462 ();
 FILLCELL_X32 FILLCELL_190_494 ();
 FILLCELL_X16 FILLCELL_190_526 ();
 FILLCELL_X8 FILLCELL_190_542 ();
 FILLCELL_X32 FILLCELL_190_552 ();
 FILLCELL_X32 FILLCELL_190_584 ();
 FILLCELL_X32 FILLCELL_190_616 ();
 FILLCELL_X32 FILLCELL_190_648 ();
 FILLCELL_X32 FILLCELL_190_680 ();
 FILLCELL_X32 FILLCELL_190_712 ();
 FILLCELL_X16 FILLCELL_190_744 ();
 FILLCELL_X8 FILLCELL_190_760 ();
 FILLCELL_X2 FILLCELL_190_768 ();
 FILLCELL_X1 FILLCELL_190_770 ();
 FILLCELL_X32 FILLCELL_190_773 ();
 FILLCELL_X32 FILLCELL_190_805 ();
 FILLCELL_X32 FILLCELL_190_837 ();
 FILLCELL_X32 FILLCELL_190_869 ();
 FILLCELL_X32 FILLCELL_190_901 ();
 FILLCELL_X32 FILLCELL_190_933 ();
 FILLCELL_X32 FILLCELL_190_965 ();
 FILLCELL_X32 FILLCELL_190_997 ();
 FILLCELL_X32 FILLCELL_190_1029 ();
 FILLCELL_X32 FILLCELL_190_1061 ();
 FILLCELL_X32 FILLCELL_190_1093 ();
 FILLCELL_X32 FILLCELL_190_1125 ();
 FILLCELL_X32 FILLCELL_190_1157 ();
 FILLCELL_X32 FILLCELL_190_1189 ();
 FILLCELL_X32 FILLCELL_190_1221 ();
 FILLCELL_X32 FILLCELL_190_1253 ();
 FILLCELL_X32 FILLCELL_190_1285 ();
 FILLCELL_X32 FILLCELL_190_1317 ();
 FILLCELL_X32 FILLCELL_190_1349 ();
 FILLCELL_X32 FILLCELL_190_1381 ();
 FILLCELL_X32 FILLCELL_190_1413 ();
 FILLCELL_X32 FILLCELL_190_1445 ();
 FILLCELL_X32 FILLCELL_190_1477 ();
 FILLCELL_X32 FILLCELL_190_1509 ();
 FILLCELL_X32 FILLCELL_190_1541 ();
 FILLCELL_X32 FILLCELL_190_1573 ();
 FILLCELL_X32 FILLCELL_190_1605 ();
 FILLCELL_X32 FILLCELL_190_1637 ();
 FILLCELL_X32 FILLCELL_190_1669 ();
 FILLCELL_X32 FILLCELL_190_1701 ();
 FILLCELL_X32 FILLCELL_190_1733 ();
 FILLCELL_X32 FILLCELL_190_1765 ();
 FILLCELL_X32 FILLCELL_190_1797 ();
 FILLCELL_X32 FILLCELL_190_1829 ();
 FILLCELL_X32 FILLCELL_190_1861 ();
 FILLCELL_X4 FILLCELL_190_1893 ();
 FILLCELL_X32 FILLCELL_191_0 ();
 FILLCELL_X32 FILLCELL_191_32 ();
 FILLCELL_X32 FILLCELL_191_64 ();
 FILLCELL_X32 FILLCELL_191_96 ();
 FILLCELL_X32 FILLCELL_191_128 ();
 FILLCELL_X32 FILLCELL_191_160 ();
 FILLCELL_X32 FILLCELL_191_192 ();
 FILLCELL_X32 FILLCELL_191_224 ();
 FILLCELL_X32 FILLCELL_191_256 ();
 FILLCELL_X32 FILLCELL_191_288 ();
 FILLCELL_X32 FILLCELL_191_320 ();
 FILLCELL_X32 FILLCELL_191_352 ();
 FILLCELL_X32 FILLCELL_191_384 ();
 FILLCELL_X32 FILLCELL_191_416 ();
 FILLCELL_X32 FILLCELL_191_448 ();
 FILLCELL_X32 FILLCELL_191_480 ();
 FILLCELL_X32 FILLCELL_191_512 ();
 FILLCELL_X32 FILLCELL_191_544 ();
 FILLCELL_X32 FILLCELL_191_576 ();
 FILLCELL_X32 FILLCELL_191_608 ();
 FILLCELL_X32 FILLCELL_191_640 ();
 FILLCELL_X32 FILLCELL_191_672 ();
 FILLCELL_X32 FILLCELL_191_704 ();
 FILLCELL_X32 FILLCELL_191_736 ();
 FILLCELL_X32 FILLCELL_191_768 ();
 FILLCELL_X32 FILLCELL_191_800 ();
 FILLCELL_X32 FILLCELL_191_832 ();
 FILLCELL_X32 FILLCELL_191_864 ();
 FILLCELL_X32 FILLCELL_191_896 ();
 FILLCELL_X32 FILLCELL_191_928 ();
 FILLCELL_X32 FILLCELL_191_960 ();
 FILLCELL_X32 FILLCELL_191_992 ();
 FILLCELL_X32 FILLCELL_191_1024 ();
 FILLCELL_X32 FILLCELL_191_1056 ();
 FILLCELL_X32 FILLCELL_191_1088 ();
 FILLCELL_X32 FILLCELL_191_1120 ();
 FILLCELL_X32 FILLCELL_191_1152 ();
 FILLCELL_X32 FILLCELL_191_1184 ();
 FILLCELL_X32 FILLCELL_191_1216 ();
 FILLCELL_X32 FILLCELL_191_1248 ();
 FILLCELL_X32 FILLCELL_191_1280 ();
 FILLCELL_X32 FILLCELL_191_1312 ();
 FILLCELL_X32 FILLCELL_191_1344 ();
 FILLCELL_X32 FILLCELL_191_1376 ();
 FILLCELL_X32 FILLCELL_191_1408 ();
 FILLCELL_X32 FILLCELL_191_1440 ();
 FILLCELL_X32 FILLCELL_191_1472 ();
 FILLCELL_X32 FILLCELL_191_1504 ();
 FILLCELL_X32 FILLCELL_191_1536 ();
 FILLCELL_X32 FILLCELL_191_1568 ();
 FILLCELL_X32 FILLCELL_191_1600 ();
 FILLCELL_X32 FILLCELL_191_1632 ();
 FILLCELL_X32 FILLCELL_191_1664 ();
 FILLCELL_X32 FILLCELL_191_1696 ();
 FILLCELL_X32 FILLCELL_191_1728 ();
 FILLCELL_X32 FILLCELL_191_1760 ();
 FILLCELL_X32 FILLCELL_191_1792 ();
 FILLCELL_X32 FILLCELL_191_1824 ();
 FILLCELL_X32 FILLCELL_191_1856 ();
 FILLCELL_X8 FILLCELL_191_1888 ();
 FILLCELL_X1 FILLCELL_191_1896 ();
 FILLCELL_X32 FILLCELL_192_0 ();
 FILLCELL_X32 FILLCELL_192_32 ();
 FILLCELL_X32 FILLCELL_192_64 ();
 FILLCELL_X32 FILLCELL_192_96 ();
 FILLCELL_X32 FILLCELL_192_128 ();
 FILLCELL_X32 FILLCELL_192_160 ();
 FILLCELL_X32 FILLCELL_192_192 ();
 FILLCELL_X32 FILLCELL_192_224 ();
 FILLCELL_X32 FILLCELL_192_256 ();
 FILLCELL_X32 FILLCELL_192_288 ();
 FILLCELL_X32 FILLCELL_192_320 ();
 FILLCELL_X32 FILLCELL_192_352 ();
 FILLCELL_X32 FILLCELL_192_384 ();
 FILLCELL_X32 FILLCELL_192_416 ();
 FILLCELL_X4 FILLCELL_192_448 ();
 FILLCELL_X32 FILLCELL_192_455 ();
 FILLCELL_X32 FILLCELL_192_487 ();
 FILLCELL_X32 FILLCELL_192_519 ();
 FILLCELL_X16 FILLCELL_192_551 ();
 FILLCELL_X2 FILLCELL_192_567 ();
 FILLCELL_X32 FILLCELL_192_574 ();
 FILLCELL_X32 FILLCELL_192_606 ();
 FILLCELL_X32 FILLCELL_192_638 ();
 FILLCELL_X32 FILLCELL_192_670 ();
 FILLCELL_X32 FILLCELL_192_702 ();
 FILLCELL_X32 FILLCELL_192_734 ();
 FILLCELL_X32 FILLCELL_192_766 ();
 FILLCELL_X32 FILLCELL_192_798 ();
 FILLCELL_X32 FILLCELL_192_830 ();
 FILLCELL_X32 FILLCELL_192_862 ();
 FILLCELL_X32 FILLCELL_192_894 ();
 FILLCELL_X32 FILLCELL_192_926 ();
 FILLCELL_X8 FILLCELL_192_958 ();
 FILLCELL_X4 FILLCELL_192_966 ();
 FILLCELL_X2 FILLCELL_192_970 ();
 FILLCELL_X32 FILLCELL_192_989 ();
 FILLCELL_X32 FILLCELL_192_1021 ();
 FILLCELL_X32 FILLCELL_192_1053 ();
 FILLCELL_X32 FILLCELL_192_1085 ();
 FILLCELL_X32 FILLCELL_192_1117 ();
 FILLCELL_X32 FILLCELL_192_1149 ();
 FILLCELL_X32 FILLCELL_192_1181 ();
 FILLCELL_X32 FILLCELL_192_1213 ();
 FILLCELL_X32 FILLCELL_192_1245 ();
 FILLCELL_X32 FILLCELL_192_1277 ();
 FILLCELL_X32 FILLCELL_192_1309 ();
 FILLCELL_X32 FILLCELL_192_1341 ();
 FILLCELL_X32 FILLCELL_192_1373 ();
 FILLCELL_X32 FILLCELL_192_1405 ();
 FILLCELL_X32 FILLCELL_192_1437 ();
 FILLCELL_X32 FILLCELL_192_1469 ();
 FILLCELL_X32 FILLCELL_192_1501 ();
 FILLCELL_X32 FILLCELL_192_1533 ();
 FILLCELL_X32 FILLCELL_192_1565 ();
 FILLCELL_X32 FILLCELL_192_1597 ();
 FILLCELL_X32 FILLCELL_192_1629 ();
 FILLCELL_X32 FILLCELL_192_1661 ();
 FILLCELL_X32 FILLCELL_192_1693 ();
 FILLCELL_X32 FILLCELL_192_1725 ();
 FILLCELL_X32 FILLCELL_192_1757 ();
 FILLCELL_X32 FILLCELL_192_1789 ();
 FILLCELL_X32 FILLCELL_192_1821 ();
 FILLCELL_X32 FILLCELL_192_1853 ();
 FILLCELL_X8 FILLCELL_192_1885 ();
 FILLCELL_X4 FILLCELL_192_1893 ();
 FILLCELL_X32 FILLCELL_193_0 ();
 FILLCELL_X32 FILLCELL_193_32 ();
 FILLCELL_X32 FILLCELL_193_64 ();
 FILLCELL_X32 FILLCELL_193_96 ();
 FILLCELL_X32 FILLCELL_193_128 ();
 FILLCELL_X32 FILLCELL_193_160 ();
 FILLCELL_X32 FILLCELL_193_192 ();
 FILLCELL_X32 FILLCELL_193_224 ();
 FILLCELL_X32 FILLCELL_193_256 ();
 FILLCELL_X32 FILLCELL_193_288 ();
 FILLCELL_X32 FILLCELL_193_320 ();
 FILLCELL_X32 FILLCELL_193_352 ();
 FILLCELL_X32 FILLCELL_193_384 ();
 FILLCELL_X32 FILLCELL_193_416 ();
 FILLCELL_X32 FILLCELL_193_448 ();
 FILLCELL_X32 FILLCELL_193_480 ();
 FILLCELL_X32 FILLCELL_193_512 ();
 FILLCELL_X32 FILLCELL_193_544 ();
 FILLCELL_X32 FILLCELL_193_576 ();
 FILLCELL_X32 FILLCELL_193_608 ();
 FILLCELL_X32 FILLCELL_193_640 ();
 FILLCELL_X32 FILLCELL_193_672 ();
 FILLCELL_X32 FILLCELL_193_704 ();
 FILLCELL_X8 FILLCELL_193_736 ();
 FILLCELL_X1 FILLCELL_193_744 ();
 FILLCELL_X32 FILLCELL_193_750 ();
 FILLCELL_X32 FILLCELL_193_782 ();
 FILLCELL_X32 FILLCELL_193_814 ();
 FILLCELL_X32 FILLCELL_193_846 ();
 FILLCELL_X32 FILLCELL_193_878 ();
 FILLCELL_X32 FILLCELL_193_910 ();
 FILLCELL_X32 FILLCELL_193_942 ();
 FILLCELL_X32 FILLCELL_193_974 ();
 FILLCELL_X32 FILLCELL_193_1006 ();
 FILLCELL_X8 FILLCELL_193_1038 ();
 FILLCELL_X2 FILLCELL_193_1046 ();
 FILLCELL_X1 FILLCELL_193_1048 ();
 FILLCELL_X32 FILLCELL_193_1062 ();
 FILLCELL_X32 FILLCELL_193_1094 ();
 FILLCELL_X32 FILLCELL_193_1126 ();
 FILLCELL_X32 FILLCELL_193_1158 ();
 FILLCELL_X32 FILLCELL_193_1190 ();
 FILLCELL_X32 FILLCELL_193_1222 ();
 FILLCELL_X32 FILLCELL_193_1254 ();
 FILLCELL_X32 FILLCELL_193_1286 ();
 FILLCELL_X32 FILLCELL_193_1318 ();
 FILLCELL_X32 FILLCELL_193_1350 ();
 FILLCELL_X32 FILLCELL_193_1382 ();
 FILLCELL_X32 FILLCELL_193_1414 ();
 FILLCELL_X32 FILLCELL_193_1446 ();
 FILLCELL_X32 FILLCELL_193_1478 ();
 FILLCELL_X32 FILLCELL_193_1510 ();
 FILLCELL_X32 FILLCELL_193_1542 ();
 FILLCELL_X32 FILLCELL_193_1574 ();
 FILLCELL_X32 FILLCELL_193_1606 ();
 FILLCELL_X32 FILLCELL_193_1638 ();
 FILLCELL_X32 FILLCELL_193_1670 ();
 FILLCELL_X32 FILLCELL_193_1702 ();
 FILLCELL_X32 FILLCELL_193_1734 ();
 FILLCELL_X32 FILLCELL_193_1766 ();
 FILLCELL_X32 FILLCELL_193_1798 ();
 FILLCELL_X32 FILLCELL_193_1830 ();
 FILLCELL_X32 FILLCELL_193_1862 ();
 FILLCELL_X2 FILLCELL_193_1894 ();
 FILLCELL_X1 FILLCELL_193_1896 ();
 FILLCELL_X32 FILLCELL_194_0 ();
 FILLCELL_X32 FILLCELL_194_32 ();
 FILLCELL_X32 FILLCELL_194_64 ();
 FILLCELL_X32 FILLCELL_194_96 ();
 FILLCELL_X32 FILLCELL_194_128 ();
 FILLCELL_X32 FILLCELL_194_160 ();
 FILLCELL_X32 FILLCELL_194_192 ();
 FILLCELL_X32 FILLCELL_194_224 ();
 FILLCELL_X32 FILLCELL_194_256 ();
 FILLCELL_X32 FILLCELL_194_288 ();
 FILLCELL_X32 FILLCELL_194_320 ();
 FILLCELL_X32 FILLCELL_194_352 ();
 FILLCELL_X32 FILLCELL_194_384 ();
 FILLCELL_X32 FILLCELL_194_416 ();
 FILLCELL_X8 FILLCELL_194_448 ();
 FILLCELL_X4 FILLCELL_194_456 ();
 FILLCELL_X32 FILLCELL_194_463 ();
 FILLCELL_X32 FILLCELL_194_495 ();
 FILLCELL_X32 FILLCELL_194_527 ();
 FILLCELL_X8 FILLCELL_194_559 ();
 FILLCELL_X4 FILLCELL_194_567 ();
 FILLCELL_X1 FILLCELL_194_571 ();
 FILLCELL_X32 FILLCELL_194_575 ();
 FILLCELL_X32 FILLCELL_194_607 ();
 FILLCELL_X32 FILLCELL_194_639 ();
 FILLCELL_X32 FILLCELL_194_671 ();
 FILLCELL_X32 FILLCELL_194_703 ();
 FILLCELL_X32 FILLCELL_194_735 ();
 FILLCELL_X32 FILLCELL_194_767 ();
 FILLCELL_X32 FILLCELL_194_799 ();
 FILLCELL_X32 FILLCELL_194_831 ();
 FILLCELL_X32 FILLCELL_194_863 ();
 FILLCELL_X32 FILLCELL_194_895 ();
 FILLCELL_X32 FILLCELL_194_927 ();
 FILLCELL_X32 FILLCELL_194_959 ();
 FILLCELL_X32 FILLCELL_194_991 ();
 FILLCELL_X32 FILLCELL_194_1023 ();
 FILLCELL_X32 FILLCELL_194_1055 ();
 FILLCELL_X16 FILLCELL_194_1087 ();
 FILLCELL_X4 FILLCELL_194_1103 ();
 FILLCELL_X32 FILLCELL_194_1120 ();
 FILLCELL_X32 FILLCELL_194_1152 ();
 FILLCELL_X32 FILLCELL_194_1184 ();
 FILLCELL_X32 FILLCELL_194_1216 ();
 FILLCELL_X32 FILLCELL_194_1248 ();
 FILLCELL_X32 FILLCELL_194_1280 ();
 FILLCELL_X32 FILLCELL_194_1312 ();
 FILLCELL_X32 FILLCELL_194_1344 ();
 FILLCELL_X32 FILLCELL_194_1376 ();
 FILLCELL_X32 FILLCELL_194_1408 ();
 FILLCELL_X32 FILLCELL_194_1440 ();
 FILLCELL_X32 FILLCELL_194_1472 ();
 FILLCELL_X32 FILLCELL_194_1504 ();
 FILLCELL_X32 FILLCELL_194_1536 ();
 FILLCELL_X32 FILLCELL_194_1568 ();
 FILLCELL_X32 FILLCELL_194_1600 ();
 FILLCELL_X32 FILLCELL_194_1632 ();
 FILLCELL_X32 FILLCELL_194_1664 ();
 FILLCELL_X32 FILLCELL_194_1696 ();
 FILLCELL_X32 FILLCELL_194_1728 ();
 FILLCELL_X32 FILLCELL_194_1760 ();
 FILLCELL_X32 FILLCELL_194_1792 ();
 FILLCELL_X32 FILLCELL_194_1824 ();
 FILLCELL_X32 FILLCELL_194_1856 ();
 FILLCELL_X8 FILLCELL_194_1888 ();
 FILLCELL_X1 FILLCELL_194_1896 ();
 FILLCELL_X32 FILLCELL_195_0 ();
 FILLCELL_X32 FILLCELL_195_32 ();
 FILLCELL_X32 FILLCELL_195_64 ();
 FILLCELL_X32 FILLCELL_195_96 ();
 FILLCELL_X32 FILLCELL_195_128 ();
 FILLCELL_X32 FILLCELL_195_160 ();
 FILLCELL_X32 FILLCELL_195_192 ();
 FILLCELL_X32 FILLCELL_195_224 ();
 FILLCELL_X32 FILLCELL_195_256 ();
 FILLCELL_X32 FILLCELL_195_288 ();
 FILLCELL_X32 FILLCELL_195_320 ();
 FILLCELL_X32 FILLCELL_195_352 ();
 FILLCELL_X32 FILLCELL_195_384 ();
 FILLCELL_X32 FILLCELL_195_416 ();
 FILLCELL_X32 FILLCELL_195_448 ();
 FILLCELL_X32 FILLCELL_195_480 ();
 FILLCELL_X32 FILLCELL_195_512 ();
 FILLCELL_X32 FILLCELL_195_544 ();
 FILLCELL_X32 FILLCELL_195_576 ();
 FILLCELL_X32 FILLCELL_195_608 ();
 FILLCELL_X8 FILLCELL_195_640 ();
 FILLCELL_X4 FILLCELL_195_648 ();
 FILLCELL_X2 FILLCELL_195_652 ();
 FILLCELL_X32 FILLCELL_195_663 ();
 FILLCELL_X32 FILLCELL_195_695 ();
 FILLCELL_X32 FILLCELL_195_727 ();
 FILLCELL_X32 FILLCELL_195_759 ();
 FILLCELL_X32 FILLCELL_195_791 ();
 FILLCELL_X32 FILLCELL_195_823 ();
 FILLCELL_X32 FILLCELL_195_855 ();
 FILLCELL_X32 FILLCELL_195_887 ();
 FILLCELL_X32 FILLCELL_195_919 ();
 FILLCELL_X32 FILLCELL_195_951 ();
 FILLCELL_X32 FILLCELL_195_983 ();
 FILLCELL_X32 FILLCELL_195_1015 ();
 FILLCELL_X32 FILLCELL_195_1047 ();
 FILLCELL_X32 FILLCELL_195_1079 ();
 FILLCELL_X32 FILLCELL_195_1111 ();
 FILLCELL_X32 FILLCELL_195_1143 ();
 FILLCELL_X32 FILLCELL_195_1175 ();
 FILLCELL_X32 FILLCELL_195_1207 ();
 FILLCELL_X32 FILLCELL_195_1239 ();
 FILLCELL_X32 FILLCELL_195_1271 ();
 FILLCELL_X32 FILLCELL_195_1303 ();
 FILLCELL_X32 FILLCELL_195_1335 ();
 FILLCELL_X32 FILLCELL_195_1367 ();
 FILLCELL_X32 FILLCELL_195_1399 ();
 FILLCELL_X32 FILLCELL_195_1431 ();
 FILLCELL_X32 FILLCELL_195_1463 ();
 FILLCELL_X32 FILLCELL_195_1495 ();
 FILLCELL_X32 FILLCELL_195_1527 ();
 FILLCELL_X32 FILLCELL_195_1559 ();
 FILLCELL_X32 FILLCELL_195_1591 ();
 FILLCELL_X32 FILLCELL_195_1623 ();
 FILLCELL_X32 FILLCELL_195_1655 ();
 FILLCELL_X32 FILLCELL_195_1687 ();
 FILLCELL_X32 FILLCELL_195_1719 ();
 FILLCELL_X32 FILLCELL_195_1751 ();
 FILLCELL_X32 FILLCELL_195_1783 ();
 FILLCELL_X32 FILLCELL_195_1815 ();
 FILLCELL_X32 FILLCELL_195_1847 ();
 FILLCELL_X16 FILLCELL_195_1879 ();
 FILLCELL_X2 FILLCELL_195_1895 ();
 FILLCELL_X32 FILLCELL_196_0 ();
 FILLCELL_X32 FILLCELL_196_32 ();
 FILLCELL_X32 FILLCELL_196_64 ();
 FILLCELL_X32 FILLCELL_196_96 ();
 FILLCELL_X32 FILLCELL_196_128 ();
 FILLCELL_X32 FILLCELL_196_160 ();
 FILLCELL_X32 FILLCELL_196_192 ();
 FILLCELL_X32 FILLCELL_196_224 ();
 FILLCELL_X32 FILLCELL_196_256 ();
 FILLCELL_X32 FILLCELL_196_288 ();
 FILLCELL_X32 FILLCELL_196_320 ();
 FILLCELL_X16 FILLCELL_196_352 ();
 FILLCELL_X1 FILLCELL_196_368 ();
 FILLCELL_X16 FILLCELL_196_373 ();
 FILLCELL_X2 FILLCELL_196_389 ();
 FILLCELL_X32 FILLCELL_196_394 ();
 FILLCELL_X32 FILLCELL_196_426 ();
 FILLCELL_X32 FILLCELL_196_458 ();
 FILLCELL_X32 FILLCELL_196_490 ();
 FILLCELL_X32 FILLCELL_196_522 ();
 FILLCELL_X32 FILLCELL_196_554 ();
 FILLCELL_X32 FILLCELL_196_586 ();
 FILLCELL_X16 FILLCELL_196_618 ();
 FILLCELL_X8 FILLCELL_196_634 ();
 FILLCELL_X2 FILLCELL_196_642 ();
 FILLCELL_X1 FILLCELL_196_644 ();
 FILLCELL_X32 FILLCELL_196_652 ();
 FILLCELL_X32 FILLCELL_196_684 ();
 FILLCELL_X32 FILLCELL_196_716 ();
 FILLCELL_X32 FILLCELL_196_748 ();
 FILLCELL_X32 FILLCELL_196_780 ();
 FILLCELL_X32 FILLCELL_196_812 ();
 FILLCELL_X32 FILLCELL_196_844 ();
 FILLCELL_X32 FILLCELL_196_876 ();
 FILLCELL_X32 FILLCELL_196_908 ();
 FILLCELL_X32 FILLCELL_196_940 ();
 FILLCELL_X32 FILLCELL_196_972 ();
 FILLCELL_X32 FILLCELL_196_1004 ();
 FILLCELL_X32 FILLCELL_196_1036 ();
 FILLCELL_X32 FILLCELL_196_1068 ();
 FILLCELL_X32 FILLCELL_196_1100 ();
 FILLCELL_X32 FILLCELL_196_1132 ();
 FILLCELL_X32 FILLCELL_196_1164 ();
 FILLCELL_X32 FILLCELL_196_1196 ();
 FILLCELL_X32 FILLCELL_196_1228 ();
 FILLCELL_X32 FILLCELL_196_1260 ();
 FILLCELL_X32 FILLCELL_196_1292 ();
 FILLCELL_X32 FILLCELL_196_1324 ();
 FILLCELL_X32 FILLCELL_196_1356 ();
 FILLCELL_X32 FILLCELL_196_1388 ();
 FILLCELL_X32 FILLCELL_196_1420 ();
 FILLCELL_X32 FILLCELL_196_1452 ();
 FILLCELL_X32 FILLCELL_196_1484 ();
 FILLCELL_X32 FILLCELL_196_1516 ();
 FILLCELL_X32 FILLCELL_196_1548 ();
 FILLCELL_X32 FILLCELL_196_1580 ();
 FILLCELL_X32 FILLCELL_196_1612 ();
 FILLCELL_X32 FILLCELL_196_1644 ();
 FILLCELL_X32 FILLCELL_196_1676 ();
 FILLCELL_X32 FILLCELL_196_1708 ();
 FILLCELL_X32 FILLCELL_196_1740 ();
 FILLCELL_X32 FILLCELL_196_1772 ();
 FILLCELL_X32 FILLCELL_196_1804 ();
 FILLCELL_X32 FILLCELL_196_1836 ();
 FILLCELL_X16 FILLCELL_196_1868 ();
 FILLCELL_X8 FILLCELL_196_1884 ();
 FILLCELL_X4 FILLCELL_196_1892 ();
 FILLCELL_X1 FILLCELL_196_1896 ();
 FILLCELL_X32 FILLCELL_197_0 ();
 FILLCELL_X32 FILLCELL_197_32 ();
 FILLCELL_X32 FILLCELL_197_64 ();
 FILLCELL_X32 FILLCELL_197_96 ();
 FILLCELL_X32 FILLCELL_197_128 ();
 FILLCELL_X32 FILLCELL_197_160 ();
 FILLCELL_X32 FILLCELL_197_192 ();
 FILLCELL_X32 FILLCELL_197_224 ();
 FILLCELL_X32 FILLCELL_197_256 ();
 FILLCELL_X32 FILLCELL_197_288 ();
 FILLCELL_X32 FILLCELL_197_320 ();
 FILLCELL_X32 FILLCELL_197_352 ();
 FILLCELL_X32 FILLCELL_197_384 ();
 FILLCELL_X16 FILLCELL_197_416 ();
 FILLCELL_X8 FILLCELL_197_432 ();
 FILLCELL_X4 FILLCELL_197_440 ();
 FILLCELL_X1 FILLCELL_197_444 ();
 FILLCELL_X32 FILLCELL_197_452 ();
 FILLCELL_X32 FILLCELL_197_484 ();
 FILLCELL_X32 FILLCELL_197_516 ();
 FILLCELL_X32 FILLCELL_197_548 ();
 FILLCELL_X32 FILLCELL_197_580 ();
 FILLCELL_X32 FILLCELL_197_612 ();
 FILLCELL_X32 FILLCELL_197_644 ();
 FILLCELL_X32 FILLCELL_197_676 ();
 FILLCELL_X32 FILLCELL_197_708 ();
 FILLCELL_X16 FILLCELL_197_740 ();
 FILLCELL_X4 FILLCELL_197_756 ();
 FILLCELL_X1 FILLCELL_197_760 ();
 FILLCELL_X32 FILLCELL_197_764 ();
 FILLCELL_X32 FILLCELL_197_796 ();
 FILLCELL_X16 FILLCELL_197_828 ();
 FILLCELL_X8 FILLCELL_197_844 ();
 FILLCELL_X4 FILLCELL_197_852 ();
 FILLCELL_X1 FILLCELL_197_856 ();
 FILLCELL_X32 FILLCELL_197_861 ();
 FILLCELL_X32 FILLCELL_197_893 ();
 FILLCELL_X32 FILLCELL_197_925 ();
 FILLCELL_X32 FILLCELL_197_957 ();
 FILLCELL_X32 FILLCELL_197_989 ();
 FILLCELL_X32 FILLCELL_197_1021 ();
 FILLCELL_X32 FILLCELL_197_1053 ();
 FILLCELL_X32 FILLCELL_197_1085 ();
 FILLCELL_X32 FILLCELL_197_1117 ();
 FILLCELL_X32 FILLCELL_197_1149 ();
 FILLCELL_X32 FILLCELL_197_1181 ();
 FILLCELL_X32 FILLCELL_197_1213 ();
 FILLCELL_X32 FILLCELL_197_1245 ();
 FILLCELL_X32 FILLCELL_197_1277 ();
 FILLCELL_X32 FILLCELL_197_1309 ();
 FILLCELL_X32 FILLCELL_197_1341 ();
 FILLCELL_X32 FILLCELL_197_1373 ();
 FILLCELL_X32 FILLCELL_197_1405 ();
 FILLCELL_X32 FILLCELL_197_1437 ();
 FILLCELL_X32 FILLCELL_197_1469 ();
 FILLCELL_X32 FILLCELL_197_1501 ();
 FILLCELL_X32 FILLCELL_197_1533 ();
 FILLCELL_X32 FILLCELL_197_1565 ();
 FILLCELL_X32 FILLCELL_197_1597 ();
 FILLCELL_X32 FILLCELL_197_1629 ();
 FILLCELL_X32 FILLCELL_197_1661 ();
 FILLCELL_X32 FILLCELL_197_1693 ();
 FILLCELL_X32 FILLCELL_197_1725 ();
 FILLCELL_X32 FILLCELL_197_1757 ();
 FILLCELL_X32 FILLCELL_197_1789 ();
 FILLCELL_X32 FILLCELL_197_1821 ();
 FILLCELL_X32 FILLCELL_197_1853 ();
 FILLCELL_X8 FILLCELL_197_1885 ();
 FILLCELL_X4 FILLCELL_197_1893 ();
 FILLCELL_X32 FILLCELL_198_0 ();
 FILLCELL_X32 FILLCELL_198_32 ();
 FILLCELL_X32 FILLCELL_198_64 ();
 FILLCELL_X32 FILLCELL_198_96 ();
 FILLCELL_X32 FILLCELL_198_128 ();
 FILLCELL_X32 FILLCELL_198_160 ();
 FILLCELL_X32 FILLCELL_198_192 ();
 FILLCELL_X32 FILLCELL_198_224 ();
 FILLCELL_X32 FILLCELL_198_256 ();
 FILLCELL_X32 FILLCELL_198_288 ();
 FILLCELL_X32 FILLCELL_198_320 ();
 FILLCELL_X32 FILLCELL_198_352 ();
 FILLCELL_X32 FILLCELL_198_384 ();
 FILLCELL_X32 FILLCELL_198_416 ();
 FILLCELL_X32 FILLCELL_198_448 ();
 FILLCELL_X32 FILLCELL_198_480 ();
 FILLCELL_X32 FILLCELL_198_512 ();
 FILLCELL_X32 FILLCELL_198_544 ();
 FILLCELL_X32 FILLCELL_198_576 ();
 FILLCELL_X32 FILLCELL_198_608 ();
 FILLCELL_X32 FILLCELL_198_640 ();
 FILLCELL_X32 FILLCELL_198_672 ();
 FILLCELL_X32 FILLCELL_198_704 ();
 FILLCELL_X32 FILLCELL_198_736 ();
 FILLCELL_X8 FILLCELL_198_768 ();
 FILLCELL_X4 FILLCELL_198_776 ();
 FILLCELL_X2 FILLCELL_198_780 ();
 FILLCELL_X32 FILLCELL_198_789 ();
 FILLCELL_X16 FILLCELL_198_821 ();
 FILLCELL_X4 FILLCELL_198_837 ();
 FILLCELL_X2 FILLCELL_198_841 ();
 FILLCELL_X32 FILLCELL_198_848 ();
 FILLCELL_X32 FILLCELL_198_880 ();
 FILLCELL_X32 FILLCELL_198_912 ();
 FILLCELL_X32 FILLCELL_198_944 ();
 FILLCELL_X32 FILLCELL_198_976 ();
 FILLCELL_X32 FILLCELL_198_1008 ();
 FILLCELL_X32 FILLCELL_198_1040 ();
 FILLCELL_X32 FILLCELL_198_1072 ();
 FILLCELL_X32 FILLCELL_198_1104 ();
 FILLCELL_X32 FILLCELL_198_1136 ();
 FILLCELL_X32 FILLCELL_198_1168 ();
 FILLCELL_X32 FILLCELL_198_1200 ();
 FILLCELL_X32 FILLCELL_198_1232 ();
 FILLCELL_X32 FILLCELL_198_1264 ();
 FILLCELL_X32 FILLCELL_198_1296 ();
 FILLCELL_X32 FILLCELL_198_1328 ();
 FILLCELL_X32 FILLCELL_198_1360 ();
 FILLCELL_X32 FILLCELL_198_1392 ();
 FILLCELL_X32 FILLCELL_198_1424 ();
 FILLCELL_X32 FILLCELL_198_1456 ();
 FILLCELL_X32 FILLCELL_198_1488 ();
 FILLCELL_X32 FILLCELL_198_1520 ();
 FILLCELL_X32 FILLCELL_198_1552 ();
 FILLCELL_X32 FILLCELL_198_1584 ();
 FILLCELL_X32 FILLCELL_198_1616 ();
 FILLCELL_X32 FILLCELL_198_1648 ();
 FILLCELL_X32 FILLCELL_198_1680 ();
 FILLCELL_X32 FILLCELL_198_1712 ();
 FILLCELL_X32 FILLCELL_198_1744 ();
 FILLCELL_X32 FILLCELL_198_1776 ();
 FILLCELL_X32 FILLCELL_198_1808 ();
 FILLCELL_X32 FILLCELL_198_1840 ();
 FILLCELL_X16 FILLCELL_198_1872 ();
 FILLCELL_X8 FILLCELL_198_1888 ();
 FILLCELL_X1 FILLCELL_198_1896 ();
 FILLCELL_X32 FILLCELL_199_0 ();
 FILLCELL_X32 FILLCELL_199_32 ();
 FILLCELL_X32 FILLCELL_199_64 ();
 FILLCELL_X32 FILLCELL_199_96 ();
 FILLCELL_X32 FILLCELL_199_128 ();
 FILLCELL_X32 FILLCELL_199_160 ();
 FILLCELL_X32 FILLCELL_199_192 ();
 FILLCELL_X2 FILLCELL_199_224 ();
 FILLCELL_X32 FILLCELL_199_229 ();
 FILLCELL_X32 FILLCELL_199_261 ();
 FILLCELL_X32 FILLCELL_199_293 ();
 FILLCELL_X32 FILLCELL_199_325 ();
 FILLCELL_X32 FILLCELL_199_357 ();
 FILLCELL_X32 FILLCELL_199_389 ();
 FILLCELL_X32 FILLCELL_199_421 ();
 FILLCELL_X32 FILLCELL_199_453 ();
 FILLCELL_X32 FILLCELL_199_485 ();
 FILLCELL_X32 FILLCELL_199_517 ();
 FILLCELL_X8 FILLCELL_199_549 ();
 FILLCELL_X2 FILLCELL_199_557 ();
 FILLCELL_X32 FILLCELL_199_576 ();
 FILLCELL_X32 FILLCELL_199_608 ();
 FILLCELL_X32 FILLCELL_199_640 ();
 FILLCELL_X8 FILLCELL_199_672 ();
 FILLCELL_X2 FILLCELL_199_680 ();
 FILLCELL_X32 FILLCELL_199_685 ();
 FILLCELL_X32 FILLCELL_199_717 ();
 FILLCELL_X32 FILLCELL_199_749 ();
 FILLCELL_X32 FILLCELL_199_781 ();
 FILLCELL_X32 FILLCELL_199_813 ();
 FILLCELL_X32 FILLCELL_199_845 ();
 FILLCELL_X32 FILLCELL_199_877 ();
 FILLCELL_X32 FILLCELL_199_909 ();
 FILLCELL_X32 FILLCELL_199_941 ();
 FILLCELL_X32 FILLCELL_199_973 ();
 FILLCELL_X32 FILLCELL_199_1005 ();
 FILLCELL_X32 FILLCELL_199_1037 ();
 FILLCELL_X32 FILLCELL_199_1069 ();
 FILLCELL_X32 FILLCELL_199_1101 ();
 FILLCELL_X32 FILLCELL_199_1133 ();
 FILLCELL_X32 FILLCELL_199_1165 ();
 FILLCELL_X32 FILLCELL_199_1197 ();
 FILLCELL_X32 FILLCELL_199_1229 ();
 FILLCELL_X32 FILLCELL_199_1261 ();
 FILLCELL_X32 FILLCELL_199_1293 ();
 FILLCELL_X32 FILLCELL_199_1325 ();
 FILLCELL_X32 FILLCELL_199_1357 ();
 FILLCELL_X32 FILLCELL_199_1389 ();
 FILLCELL_X32 FILLCELL_199_1421 ();
 FILLCELL_X32 FILLCELL_199_1453 ();
 FILLCELL_X32 FILLCELL_199_1485 ();
 FILLCELL_X32 FILLCELL_199_1517 ();
 FILLCELL_X32 FILLCELL_199_1549 ();
 FILLCELL_X32 FILLCELL_199_1581 ();
 FILLCELL_X32 FILLCELL_199_1613 ();
 FILLCELL_X32 FILLCELL_199_1645 ();
 FILLCELL_X32 FILLCELL_199_1677 ();
 FILLCELL_X32 FILLCELL_199_1709 ();
 FILLCELL_X32 FILLCELL_199_1741 ();
 FILLCELL_X32 FILLCELL_199_1773 ();
 FILLCELL_X32 FILLCELL_199_1805 ();
 FILLCELL_X32 FILLCELL_199_1837 ();
 FILLCELL_X16 FILLCELL_199_1869 ();
 FILLCELL_X8 FILLCELL_199_1885 ();
 FILLCELL_X4 FILLCELL_199_1893 ();
 FILLCELL_X32 FILLCELL_200_0 ();
 FILLCELL_X32 FILLCELL_200_32 ();
 FILLCELL_X32 FILLCELL_200_64 ();
 FILLCELL_X32 FILLCELL_200_96 ();
 FILLCELL_X32 FILLCELL_200_128 ();
 FILLCELL_X32 FILLCELL_200_160 ();
 FILLCELL_X32 FILLCELL_200_192 ();
 FILLCELL_X32 FILLCELL_200_224 ();
 FILLCELL_X32 FILLCELL_200_256 ();
 FILLCELL_X32 FILLCELL_200_288 ();
 FILLCELL_X32 FILLCELL_200_320 ();
 FILLCELL_X32 FILLCELL_200_352 ();
 FILLCELL_X32 FILLCELL_200_384 ();
 FILLCELL_X32 FILLCELL_200_416 ();
 FILLCELL_X32 FILLCELL_200_448 ();
 FILLCELL_X32 FILLCELL_200_480 ();
 FILLCELL_X32 FILLCELL_200_512 ();
 FILLCELL_X32 FILLCELL_200_544 ();
 FILLCELL_X32 FILLCELL_200_576 ();
 FILLCELL_X32 FILLCELL_200_608 ();
 FILLCELL_X32 FILLCELL_200_640 ();
 FILLCELL_X32 FILLCELL_200_672 ();
 FILLCELL_X32 FILLCELL_200_704 ();
 FILLCELL_X32 FILLCELL_200_736 ();
 FILLCELL_X32 FILLCELL_200_768 ();
 FILLCELL_X32 FILLCELL_200_800 ();
 FILLCELL_X32 FILLCELL_200_832 ();
 FILLCELL_X32 FILLCELL_200_864 ();
 FILLCELL_X4 FILLCELL_200_896 ();
 FILLCELL_X1 FILLCELL_200_900 ();
 FILLCELL_X32 FILLCELL_200_904 ();
 FILLCELL_X32 FILLCELL_200_936 ();
 FILLCELL_X32 FILLCELL_200_968 ();
 FILLCELL_X32 FILLCELL_200_1000 ();
 FILLCELL_X32 FILLCELL_200_1032 ();
 FILLCELL_X32 FILLCELL_200_1064 ();
 FILLCELL_X32 FILLCELL_200_1096 ();
 FILLCELL_X32 FILLCELL_200_1128 ();
 FILLCELL_X32 FILLCELL_200_1160 ();
 FILLCELL_X32 FILLCELL_200_1192 ();
 FILLCELL_X32 FILLCELL_200_1224 ();
 FILLCELL_X32 FILLCELL_200_1256 ();
 FILLCELL_X32 FILLCELL_200_1288 ();
 FILLCELL_X32 FILLCELL_200_1320 ();
 FILLCELL_X32 FILLCELL_200_1352 ();
 FILLCELL_X32 FILLCELL_200_1384 ();
 FILLCELL_X32 FILLCELL_200_1416 ();
 FILLCELL_X32 FILLCELL_200_1448 ();
 FILLCELL_X32 FILLCELL_200_1480 ();
 FILLCELL_X32 FILLCELL_200_1512 ();
 FILLCELL_X32 FILLCELL_200_1544 ();
 FILLCELL_X32 FILLCELL_200_1576 ();
 FILLCELL_X32 FILLCELL_200_1608 ();
 FILLCELL_X32 FILLCELL_200_1640 ();
 FILLCELL_X32 FILLCELL_200_1672 ();
 FILLCELL_X32 FILLCELL_200_1704 ();
 FILLCELL_X32 FILLCELL_200_1736 ();
 FILLCELL_X32 FILLCELL_200_1768 ();
 FILLCELL_X32 FILLCELL_200_1800 ();
 FILLCELL_X32 FILLCELL_200_1832 ();
 FILLCELL_X32 FILLCELL_200_1864 ();
 FILLCELL_X1 FILLCELL_200_1896 ();
 FILLCELL_X32 FILLCELL_201_0 ();
 FILLCELL_X32 FILLCELL_201_32 ();
 FILLCELL_X32 FILLCELL_201_64 ();
 FILLCELL_X32 FILLCELL_201_96 ();
 FILLCELL_X32 FILLCELL_201_128 ();
 FILLCELL_X32 FILLCELL_201_160 ();
 FILLCELL_X32 FILLCELL_201_192 ();
 FILLCELL_X32 FILLCELL_201_224 ();
 FILLCELL_X32 FILLCELL_201_256 ();
 FILLCELL_X32 FILLCELL_201_288 ();
 FILLCELL_X32 FILLCELL_201_320 ();
 FILLCELL_X32 FILLCELL_201_352 ();
 FILLCELL_X32 FILLCELL_201_384 ();
 FILLCELL_X32 FILLCELL_201_416 ();
 FILLCELL_X32 FILLCELL_201_448 ();
 FILLCELL_X32 FILLCELL_201_480 ();
 FILLCELL_X32 FILLCELL_201_512 ();
 FILLCELL_X32 FILLCELL_201_544 ();
 FILLCELL_X32 FILLCELL_201_576 ();
 FILLCELL_X32 FILLCELL_201_608 ();
 FILLCELL_X32 FILLCELL_201_640 ();
 FILLCELL_X32 FILLCELL_201_672 ();
 FILLCELL_X32 FILLCELL_201_704 ();
 FILLCELL_X32 FILLCELL_201_736 ();
 FILLCELL_X32 FILLCELL_201_768 ();
 FILLCELL_X32 FILLCELL_201_800 ();
 FILLCELL_X32 FILLCELL_201_832 ();
 FILLCELL_X32 FILLCELL_201_864 ();
 FILLCELL_X32 FILLCELL_201_896 ();
 FILLCELL_X32 FILLCELL_201_928 ();
 FILLCELL_X32 FILLCELL_201_960 ();
 FILLCELL_X32 FILLCELL_201_992 ();
 FILLCELL_X32 FILLCELL_201_1024 ();
 FILLCELL_X32 FILLCELL_201_1056 ();
 FILLCELL_X32 FILLCELL_201_1088 ();
 FILLCELL_X32 FILLCELL_201_1120 ();
 FILLCELL_X32 FILLCELL_201_1152 ();
 FILLCELL_X32 FILLCELL_201_1184 ();
 FILLCELL_X32 FILLCELL_201_1216 ();
 FILLCELL_X32 FILLCELL_201_1248 ();
 FILLCELL_X32 FILLCELL_201_1280 ();
 FILLCELL_X32 FILLCELL_201_1312 ();
 FILLCELL_X32 FILLCELL_201_1344 ();
 FILLCELL_X32 FILLCELL_201_1376 ();
 FILLCELL_X32 FILLCELL_201_1408 ();
 FILLCELL_X32 FILLCELL_201_1440 ();
 FILLCELL_X32 FILLCELL_201_1472 ();
 FILLCELL_X32 FILLCELL_201_1504 ();
 FILLCELL_X32 FILLCELL_201_1536 ();
 FILLCELL_X32 FILLCELL_201_1568 ();
 FILLCELL_X32 FILLCELL_201_1600 ();
 FILLCELL_X32 FILLCELL_201_1632 ();
 FILLCELL_X32 FILLCELL_201_1664 ();
 FILLCELL_X32 FILLCELL_201_1696 ();
 FILLCELL_X32 FILLCELL_201_1728 ();
 FILLCELL_X32 FILLCELL_201_1760 ();
 FILLCELL_X32 FILLCELL_201_1792 ();
 FILLCELL_X32 FILLCELL_201_1824 ();
 FILLCELL_X32 FILLCELL_201_1856 ();
 FILLCELL_X8 FILLCELL_201_1888 ();
 FILLCELL_X1 FILLCELL_201_1896 ();
 FILLCELL_X32 FILLCELL_202_0 ();
 FILLCELL_X32 FILLCELL_202_32 ();
 FILLCELL_X32 FILLCELL_202_64 ();
 FILLCELL_X32 FILLCELL_202_96 ();
 FILLCELL_X32 FILLCELL_202_128 ();
 FILLCELL_X32 FILLCELL_202_160 ();
 FILLCELL_X32 FILLCELL_202_192 ();
 FILLCELL_X32 FILLCELL_202_224 ();
 FILLCELL_X32 FILLCELL_202_256 ();
 FILLCELL_X32 FILLCELL_202_288 ();
 FILLCELL_X32 FILLCELL_202_320 ();
 FILLCELL_X32 FILLCELL_202_352 ();
 FILLCELL_X32 FILLCELL_202_384 ();
 FILLCELL_X16 FILLCELL_202_416 ();
 FILLCELL_X8 FILLCELL_202_432 ();
 FILLCELL_X4 FILLCELL_202_440 ();
 FILLCELL_X1 FILLCELL_202_444 ();
 FILLCELL_X32 FILLCELL_202_462 ();
 FILLCELL_X32 FILLCELL_202_494 ();
 FILLCELL_X32 FILLCELL_202_526 ();
 FILLCELL_X32 FILLCELL_202_558 ();
 FILLCELL_X32 FILLCELL_202_590 ();
 FILLCELL_X32 FILLCELL_202_622 ();
 FILLCELL_X32 FILLCELL_202_654 ();
 FILLCELL_X32 FILLCELL_202_686 ();
 FILLCELL_X32 FILLCELL_202_718 ();
 FILLCELL_X8 FILLCELL_202_750 ();
 FILLCELL_X2 FILLCELL_202_758 ();
 FILLCELL_X1 FILLCELL_202_760 ();
 FILLCELL_X32 FILLCELL_202_778 ();
 FILLCELL_X32 FILLCELL_202_810 ();
 FILLCELL_X32 FILLCELL_202_842 ();
 FILLCELL_X32 FILLCELL_202_874 ();
 FILLCELL_X32 FILLCELL_202_906 ();
 FILLCELL_X32 FILLCELL_202_938 ();
 FILLCELL_X32 FILLCELL_202_970 ();
 FILLCELL_X32 FILLCELL_202_1002 ();
 FILLCELL_X32 FILLCELL_202_1034 ();
 FILLCELL_X32 FILLCELL_202_1066 ();
 FILLCELL_X32 FILLCELL_202_1098 ();
 FILLCELL_X32 FILLCELL_202_1130 ();
 FILLCELL_X32 FILLCELL_202_1162 ();
 FILLCELL_X32 FILLCELL_202_1194 ();
 FILLCELL_X32 FILLCELL_202_1226 ();
 FILLCELL_X32 FILLCELL_202_1258 ();
 FILLCELL_X32 FILLCELL_202_1290 ();
 FILLCELL_X32 FILLCELL_202_1322 ();
 FILLCELL_X32 FILLCELL_202_1354 ();
 FILLCELL_X32 FILLCELL_202_1386 ();
 FILLCELL_X32 FILLCELL_202_1418 ();
 FILLCELL_X32 FILLCELL_202_1450 ();
 FILLCELL_X32 FILLCELL_202_1482 ();
 FILLCELL_X32 FILLCELL_202_1514 ();
 FILLCELL_X32 FILLCELL_202_1546 ();
 FILLCELL_X32 FILLCELL_202_1578 ();
 FILLCELL_X32 FILLCELL_202_1610 ();
 FILLCELL_X32 FILLCELL_202_1642 ();
 FILLCELL_X32 FILLCELL_202_1674 ();
 FILLCELL_X32 FILLCELL_202_1706 ();
 FILLCELL_X32 FILLCELL_202_1738 ();
 FILLCELL_X32 FILLCELL_202_1770 ();
 FILLCELL_X32 FILLCELL_202_1802 ();
 FILLCELL_X32 FILLCELL_202_1834 ();
 FILLCELL_X16 FILLCELL_202_1866 ();
 FILLCELL_X8 FILLCELL_202_1882 ();
 FILLCELL_X4 FILLCELL_202_1890 ();
 FILLCELL_X2 FILLCELL_202_1894 ();
 FILLCELL_X1 FILLCELL_202_1896 ();
 FILLCELL_X32 FILLCELL_203_0 ();
 FILLCELL_X32 FILLCELL_203_32 ();
 FILLCELL_X32 FILLCELL_203_64 ();
 FILLCELL_X32 FILLCELL_203_96 ();
 FILLCELL_X32 FILLCELL_203_128 ();
 FILLCELL_X32 FILLCELL_203_160 ();
 FILLCELL_X32 FILLCELL_203_192 ();
 FILLCELL_X32 FILLCELL_203_224 ();
 FILLCELL_X32 FILLCELL_203_256 ();
 FILLCELL_X32 FILLCELL_203_288 ();
 FILLCELL_X32 FILLCELL_203_320 ();
 FILLCELL_X32 FILLCELL_203_352 ();
 FILLCELL_X32 FILLCELL_203_384 ();
 FILLCELL_X32 FILLCELL_203_416 ();
 FILLCELL_X32 FILLCELL_203_448 ();
 FILLCELL_X32 FILLCELL_203_480 ();
 FILLCELL_X32 FILLCELL_203_512 ();
 FILLCELL_X32 FILLCELL_203_544 ();
 FILLCELL_X32 FILLCELL_203_576 ();
 FILLCELL_X32 FILLCELL_203_608 ();
 FILLCELL_X32 FILLCELL_203_640 ();
 FILLCELL_X32 FILLCELL_203_672 ();
 FILLCELL_X32 FILLCELL_203_704 ();
 FILLCELL_X32 FILLCELL_203_736 ();
 FILLCELL_X32 FILLCELL_203_768 ();
 FILLCELL_X32 FILLCELL_203_800 ();
 FILLCELL_X32 FILLCELL_203_832 ();
 FILLCELL_X32 FILLCELL_203_864 ();
 FILLCELL_X32 FILLCELL_203_896 ();
 FILLCELL_X32 FILLCELL_203_928 ();
 FILLCELL_X32 FILLCELL_203_960 ();
 FILLCELL_X32 FILLCELL_203_992 ();
 FILLCELL_X32 FILLCELL_203_1024 ();
 FILLCELL_X32 FILLCELL_203_1056 ();
 FILLCELL_X32 FILLCELL_203_1088 ();
 FILLCELL_X32 FILLCELL_203_1120 ();
 FILLCELL_X32 FILLCELL_203_1152 ();
 FILLCELL_X32 FILLCELL_203_1184 ();
 FILLCELL_X32 FILLCELL_203_1216 ();
 FILLCELL_X32 FILLCELL_203_1248 ();
 FILLCELL_X32 FILLCELL_203_1280 ();
 FILLCELL_X32 FILLCELL_203_1312 ();
 FILLCELL_X32 FILLCELL_203_1344 ();
 FILLCELL_X32 FILLCELL_203_1376 ();
 FILLCELL_X32 FILLCELL_203_1408 ();
 FILLCELL_X32 FILLCELL_203_1440 ();
 FILLCELL_X32 FILLCELL_203_1472 ();
 FILLCELL_X32 FILLCELL_203_1504 ();
 FILLCELL_X32 FILLCELL_203_1536 ();
 FILLCELL_X32 FILLCELL_203_1568 ();
 FILLCELL_X32 FILLCELL_203_1600 ();
 FILLCELL_X32 FILLCELL_203_1632 ();
 FILLCELL_X32 FILLCELL_203_1664 ();
 FILLCELL_X32 FILLCELL_203_1696 ();
 FILLCELL_X32 FILLCELL_203_1728 ();
 FILLCELL_X32 FILLCELL_203_1760 ();
 FILLCELL_X32 FILLCELL_203_1792 ();
 FILLCELL_X32 FILLCELL_203_1824 ();
 FILLCELL_X32 FILLCELL_203_1856 ();
 FILLCELL_X8 FILLCELL_203_1888 ();
 FILLCELL_X1 FILLCELL_203_1896 ();
 FILLCELL_X32 FILLCELL_204_0 ();
 FILLCELL_X32 FILLCELL_204_32 ();
 FILLCELL_X32 FILLCELL_204_64 ();
 FILLCELL_X32 FILLCELL_204_96 ();
 FILLCELL_X32 FILLCELL_204_128 ();
 FILLCELL_X32 FILLCELL_204_160 ();
 FILLCELL_X32 FILLCELL_204_192 ();
 FILLCELL_X32 FILLCELL_204_224 ();
 FILLCELL_X32 FILLCELL_204_256 ();
 FILLCELL_X32 FILLCELL_204_288 ();
 FILLCELL_X32 FILLCELL_204_320 ();
 FILLCELL_X32 FILLCELL_204_352 ();
 FILLCELL_X32 FILLCELL_204_384 ();
 FILLCELL_X32 FILLCELL_204_416 ();
 FILLCELL_X32 FILLCELL_204_448 ();
 FILLCELL_X32 FILLCELL_204_480 ();
 FILLCELL_X32 FILLCELL_204_512 ();
 FILLCELL_X32 FILLCELL_204_544 ();
 FILLCELL_X32 FILLCELL_204_576 ();
 FILLCELL_X32 FILLCELL_204_608 ();
 FILLCELL_X32 FILLCELL_204_640 ();
 FILLCELL_X32 FILLCELL_204_672 ();
 FILLCELL_X32 FILLCELL_204_704 ();
 FILLCELL_X32 FILLCELL_204_736 ();
 FILLCELL_X32 FILLCELL_204_768 ();
 FILLCELL_X32 FILLCELL_204_800 ();
 FILLCELL_X32 FILLCELL_204_832 ();
 FILLCELL_X32 FILLCELL_204_864 ();
 FILLCELL_X32 FILLCELL_204_896 ();
 FILLCELL_X32 FILLCELL_204_928 ();
 FILLCELL_X32 FILLCELL_204_960 ();
 FILLCELL_X32 FILLCELL_204_992 ();
 FILLCELL_X32 FILLCELL_204_1024 ();
 FILLCELL_X32 FILLCELL_204_1056 ();
 FILLCELL_X32 FILLCELL_204_1088 ();
 FILLCELL_X32 FILLCELL_204_1120 ();
 FILLCELL_X32 FILLCELL_204_1152 ();
 FILLCELL_X32 FILLCELL_204_1184 ();
 FILLCELL_X32 FILLCELL_204_1216 ();
 FILLCELL_X32 FILLCELL_204_1248 ();
 FILLCELL_X32 FILLCELL_204_1280 ();
 FILLCELL_X32 FILLCELL_204_1312 ();
 FILLCELL_X32 FILLCELL_204_1344 ();
 FILLCELL_X32 FILLCELL_204_1376 ();
 FILLCELL_X32 FILLCELL_204_1408 ();
 FILLCELL_X32 FILLCELL_204_1440 ();
 FILLCELL_X32 FILLCELL_204_1472 ();
 FILLCELL_X32 FILLCELL_204_1504 ();
 FILLCELL_X32 FILLCELL_204_1536 ();
 FILLCELL_X32 FILLCELL_204_1568 ();
 FILLCELL_X32 FILLCELL_204_1600 ();
 FILLCELL_X32 FILLCELL_204_1632 ();
 FILLCELL_X32 FILLCELL_204_1664 ();
 FILLCELL_X32 FILLCELL_204_1696 ();
 FILLCELL_X32 FILLCELL_204_1728 ();
 FILLCELL_X32 FILLCELL_204_1760 ();
 FILLCELL_X32 FILLCELL_204_1792 ();
 FILLCELL_X32 FILLCELL_204_1824 ();
 FILLCELL_X32 FILLCELL_204_1856 ();
 FILLCELL_X8 FILLCELL_204_1888 ();
 FILLCELL_X1 FILLCELL_204_1896 ();
 FILLCELL_X32 FILLCELL_205_0 ();
 FILLCELL_X32 FILLCELL_205_32 ();
 FILLCELL_X32 FILLCELL_205_64 ();
 FILLCELL_X32 FILLCELL_205_96 ();
 FILLCELL_X32 FILLCELL_205_128 ();
 FILLCELL_X32 FILLCELL_205_160 ();
 FILLCELL_X32 FILLCELL_205_192 ();
 FILLCELL_X32 FILLCELL_205_224 ();
 FILLCELL_X32 FILLCELL_205_256 ();
 FILLCELL_X32 FILLCELL_205_288 ();
 FILLCELL_X32 FILLCELL_205_320 ();
 FILLCELL_X32 FILLCELL_205_352 ();
 FILLCELL_X32 FILLCELL_205_384 ();
 FILLCELL_X32 FILLCELL_205_416 ();
 FILLCELL_X32 FILLCELL_205_448 ();
 FILLCELL_X32 FILLCELL_205_480 ();
 FILLCELL_X32 FILLCELL_205_512 ();
 FILLCELL_X32 FILLCELL_205_544 ();
 FILLCELL_X32 FILLCELL_205_576 ();
 FILLCELL_X32 FILLCELL_205_608 ();
 FILLCELL_X32 FILLCELL_205_640 ();
 FILLCELL_X32 FILLCELL_205_672 ();
 FILLCELL_X32 FILLCELL_205_704 ();
 FILLCELL_X32 FILLCELL_205_736 ();
 FILLCELL_X32 FILLCELL_205_768 ();
 FILLCELL_X32 FILLCELL_205_800 ();
 FILLCELL_X32 FILLCELL_205_832 ();
 FILLCELL_X32 FILLCELL_205_864 ();
 FILLCELL_X32 FILLCELL_205_896 ();
 FILLCELL_X32 FILLCELL_205_928 ();
 FILLCELL_X32 FILLCELL_205_960 ();
 FILLCELL_X32 FILLCELL_205_992 ();
 FILLCELL_X32 FILLCELL_205_1024 ();
 FILLCELL_X32 FILLCELL_205_1056 ();
 FILLCELL_X32 FILLCELL_205_1088 ();
 FILLCELL_X32 FILLCELL_205_1120 ();
 FILLCELL_X32 FILLCELL_205_1152 ();
 FILLCELL_X32 FILLCELL_205_1184 ();
 FILLCELL_X32 FILLCELL_205_1216 ();
 FILLCELL_X32 FILLCELL_205_1248 ();
 FILLCELL_X32 FILLCELL_205_1280 ();
 FILLCELL_X32 FILLCELL_205_1312 ();
 FILLCELL_X32 FILLCELL_205_1344 ();
 FILLCELL_X32 FILLCELL_205_1376 ();
 FILLCELL_X32 FILLCELL_205_1408 ();
 FILLCELL_X32 FILLCELL_205_1440 ();
 FILLCELL_X32 FILLCELL_205_1472 ();
 FILLCELL_X32 FILLCELL_205_1504 ();
 FILLCELL_X32 FILLCELL_205_1536 ();
 FILLCELL_X32 FILLCELL_205_1568 ();
 FILLCELL_X32 FILLCELL_205_1600 ();
 FILLCELL_X32 FILLCELL_205_1632 ();
 FILLCELL_X32 FILLCELL_205_1664 ();
 FILLCELL_X32 FILLCELL_205_1696 ();
 FILLCELL_X32 FILLCELL_205_1728 ();
 FILLCELL_X32 FILLCELL_205_1760 ();
 FILLCELL_X32 FILLCELL_205_1792 ();
 FILLCELL_X32 FILLCELL_205_1824 ();
 FILLCELL_X32 FILLCELL_205_1856 ();
 FILLCELL_X8 FILLCELL_205_1888 ();
 FILLCELL_X1 FILLCELL_205_1896 ();
 FILLCELL_X32 FILLCELL_206_0 ();
 FILLCELL_X32 FILLCELL_206_32 ();
 FILLCELL_X32 FILLCELL_206_64 ();
 FILLCELL_X32 FILLCELL_206_96 ();
 FILLCELL_X32 FILLCELL_206_128 ();
 FILLCELL_X32 FILLCELL_206_160 ();
 FILLCELL_X32 FILLCELL_206_192 ();
 FILLCELL_X32 FILLCELL_206_224 ();
 FILLCELL_X32 FILLCELL_206_256 ();
 FILLCELL_X32 FILLCELL_206_288 ();
 FILLCELL_X32 FILLCELL_206_320 ();
 FILLCELL_X32 FILLCELL_206_352 ();
 FILLCELL_X32 FILLCELL_206_384 ();
 FILLCELL_X32 FILLCELL_206_416 ();
 FILLCELL_X32 FILLCELL_206_448 ();
 FILLCELL_X32 FILLCELL_206_480 ();
 FILLCELL_X32 FILLCELL_206_512 ();
 FILLCELL_X32 FILLCELL_206_544 ();
 FILLCELL_X32 FILLCELL_206_576 ();
 FILLCELL_X32 FILLCELL_206_608 ();
 FILLCELL_X32 FILLCELL_206_640 ();
 FILLCELL_X32 FILLCELL_206_672 ();
 FILLCELL_X32 FILLCELL_206_704 ();
 FILLCELL_X32 FILLCELL_206_736 ();
 FILLCELL_X32 FILLCELL_206_768 ();
 FILLCELL_X32 FILLCELL_206_800 ();
 FILLCELL_X32 FILLCELL_206_832 ();
 FILLCELL_X32 FILLCELL_206_864 ();
 FILLCELL_X32 FILLCELL_206_896 ();
 FILLCELL_X32 FILLCELL_206_928 ();
 FILLCELL_X32 FILLCELL_206_960 ();
 FILLCELL_X32 FILLCELL_206_992 ();
 FILLCELL_X32 FILLCELL_206_1024 ();
 FILLCELL_X32 FILLCELL_206_1056 ();
 FILLCELL_X32 FILLCELL_206_1088 ();
 FILLCELL_X32 FILLCELL_206_1120 ();
 FILLCELL_X32 FILLCELL_206_1152 ();
 FILLCELL_X32 FILLCELL_206_1184 ();
 FILLCELL_X32 FILLCELL_206_1216 ();
 FILLCELL_X32 FILLCELL_206_1248 ();
 FILLCELL_X32 FILLCELL_206_1280 ();
 FILLCELL_X32 FILLCELL_206_1312 ();
 FILLCELL_X32 FILLCELL_206_1344 ();
 FILLCELL_X32 FILLCELL_206_1376 ();
 FILLCELL_X32 FILLCELL_206_1408 ();
 FILLCELL_X32 FILLCELL_206_1440 ();
 FILLCELL_X32 FILLCELL_206_1472 ();
 FILLCELL_X32 FILLCELL_206_1504 ();
 FILLCELL_X32 FILLCELL_206_1536 ();
 FILLCELL_X32 FILLCELL_206_1568 ();
 FILLCELL_X32 FILLCELL_206_1600 ();
 FILLCELL_X32 FILLCELL_206_1632 ();
 FILLCELL_X32 FILLCELL_206_1664 ();
 FILLCELL_X32 FILLCELL_206_1696 ();
 FILLCELL_X32 FILLCELL_206_1728 ();
 FILLCELL_X32 FILLCELL_206_1760 ();
 FILLCELL_X32 FILLCELL_206_1792 ();
 FILLCELL_X32 FILLCELL_206_1824 ();
 FILLCELL_X32 FILLCELL_206_1856 ();
 FILLCELL_X8 FILLCELL_206_1888 ();
 FILLCELL_X1 FILLCELL_206_1896 ();
 FILLCELL_X32 FILLCELL_207_0 ();
 FILLCELL_X32 FILLCELL_207_32 ();
 FILLCELL_X32 FILLCELL_207_64 ();
 FILLCELL_X32 FILLCELL_207_96 ();
 FILLCELL_X32 FILLCELL_207_128 ();
 FILLCELL_X32 FILLCELL_207_160 ();
 FILLCELL_X32 FILLCELL_207_192 ();
 FILLCELL_X32 FILLCELL_207_224 ();
 FILLCELL_X32 FILLCELL_207_256 ();
 FILLCELL_X32 FILLCELL_207_288 ();
 FILLCELL_X32 FILLCELL_207_320 ();
 FILLCELL_X32 FILLCELL_207_352 ();
 FILLCELL_X32 FILLCELL_207_384 ();
 FILLCELL_X32 FILLCELL_207_416 ();
 FILLCELL_X32 FILLCELL_207_448 ();
 FILLCELL_X32 FILLCELL_207_480 ();
 FILLCELL_X32 FILLCELL_207_512 ();
 FILLCELL_X32 FILLCELL_207_544 ();
 FILLCELL_X32 FILLCELL_207_576 ();
 FILLCELL_X32 FILLCELL_207_608 ();
 FILLCELL_X32 FILLCELL_207_640 ();
 FILLCELL_X32 FILLCELL_207_672 ();
 FILLCELL_X32 FILLCELL_207_704 ();
 FILLCELL_X32 FILLCELL_207_736 ();
 FILLCELL_X32 FILLCELL_207_768 ();
 FILLCELL_X32 FILLCELL_207_800 ();
 FILLCELL_X32 FILLCELL_207_832 ();
 FILLCELL_X32 FILLCELL_207_864 ();
 FILLCELL_X32 FILLCELL_207_896 ();
 FILLCELL_X32 FILLCELL_207_928 ();
 FILLCELL_X32 FILLCELL_207_960 ();
 FILLCELL_X32 FILLCELL_207_992 ();
 FILLCELL_X32 FILLCELL_207_1024 ();
 FILLCELL_X32 FILLCELL_207_1056 ();
 FILLCELL_X32 FILLCELL_207_1088 ();
 FILLCELL_X32 FILLCELL_207_1120 ();
 FILLCELL_X32 FILLCELL_207_1152 ();
 FILLCELL_X32 FILLCELL_207_1184 ();
 FILLCELL_X32 FILLCELL_207_1216 ();
 FILLCELL_X32 FILLCELL_207_1248 ();
 FILLCELL_X32 FILLCELL_207_1280 ();
 FILLCELL_X32 FILLCELL_207_1312 ();
 FILLCELL_X32 FILLCELL_207_1344 ();
 FILLCELL_X32 FILLCELL_207_1376 ();
 FILLCELL_X32 FILLCELL_207_1408 ();
 FILLCELL_X32 FILLCELL_207_1440 ();
 FILLCELL_X32 FILLCELL_207_1472 ();
 FILLCELL_X32 FILLCELL_207_1504 ();
 FILLCELL_X32 FILLCELL_207_1536 ();
 FILLCELL_X32 FILLCELL_207_1568 ();
 FILLCELL_X32 FILLCELL_207_1600 ();
 FILLCELL_X32 FILLCELL_207_1632 ();
 FILLCELL_X32 FILLCELL_207_1664 ();
 FILLCELL_X32 FILLCELL_207_1696 ();
 FILLCELL_X32 FILLCELL_207_1728 ();
 FILLCELL_X32 FILLCELL_207_1760 ();
 FILLCELL_X32 FILLCELL_207_1792 ();
 FILLCELL_X32 FILLCELL_207_1824 ();
 FILLCELL_X32 FILLCELL_207_1856 ();
 FILLCELL_X8 FILLCELL_207_1888 ();
 FILLCELL_X1 FILLCELL_207_1896 ();
 FILLCELL_X32 FILLCELL_208_0 ();
 FILLCELL_X32 FILLCELL_208_32 ();
 FILLCELL_X32 FILLCELL_208_64 ();
 FILLCELL_X32 FILLCELL_208_96 ();
 FILLCELL_X32 FILLCELL_208_128 ();
 FILLCELL_X32 FILLCELL_208_160 ();
 FILLCELL_X32 FILLCELL_208_192 ();
 FILLCELL_X32 FILLCELL_208_224 ();
 FILLCELL_X32 FILLCELL_208_256 ();
 FILLCELL_X32 FILLCELL_208_288 ();
 FILLCELL_X32 FILLCELL_208_320 ();
 FILLCELL_X32 FILLCELL_208_352 ();
 FILLCELL_X32 FILLCELL_208_384 ();
 FILLCELL_X32 FILLCELL_208_416 ();
 FILLCELL_X32 FILLCELL_208_448 ();
 FILLCELL_X32 FILLCELL_208_480 ();
 FILLCELL_X32 FILLCELL_208_512 ();
 FILLCELL_X32 FILLCELL_208_544 ();
 FILLCELL_X32 FILLCELL_208_576 ();
 FILLCELL_X32 FILLCELL_208_608 ();
 FILLCELL_X32 FILLCELL_208_640 ();
 FILLCELL_X32 FILLCELL_208_672 ();
 FILLCELL_X32 FILLCELL_208_704 ();
 FILLCELL_X32 FILLCELL_208_736 ();
 FILLCELL_X32 FILLCELL_208_768 ();
 FILLCELL_X32 FILLCELL_208_800 ();
 FILLCELL_X32 FILLCELL_208_832 ();
 FILLCELL_X32 FILLCELL_208_864 ();
 FILLCELL_X32 FILLCELL_208_896 ();
 FILLCELL_X32 FILLCELL_208_928 ();
 FILLCELL_X32 FILLCELL_208_960 ();
 FILLCELL_X32 FILLCELL_208_992 ();
 FILLCELL_X32 FILLCELL_208_1024 ();
 FILLCELL_X32 FILLCELL_208_1056 ();
 FILLCELL_X32 FILLCELL_208_1088 ();
 FILLCELL_X32 FILLCELL_208_1120 ();
 FILLCELL_X32 FILLCELL_208_1152 ();
 FILLCELL_X32 FILLCELL_208_1184 ();
 FILLCELL_X32 FILLCELL_208_1216 ();
 FILLCELL_X32 FILLCELL_208_1248 ();
 FILLCELL_X32 FILLCELL_208_1280 ();
 FILLCELL_X32 FILLCELL_208_1312 ();
 FILLCELL_X32 FILLCELL_208_1344 ();
 FILLCELL_X32 FILLCELL_208_1376 ();
 FILLCELL_X32 FILLCELL_208_1408 ();
 FILLCELL_X32 FILLCELL_208_1440 ();
 FILLCELL_X32 FILLCELL_208_1472 ();
 FILLCELL_X32 FILLCELL_208_1504 ();
 FILLCELL_X32 FILLCELL_208_1536 ();
 FILLCELL_X32 FILLCELL_208_1568 ();
 FILLCELL_X32 FILLCELL_208_1600 ();
 FILLCELL_X32 FILLCELL_208_1632 ();
 FILLCELL_X32 FILLCELL_208_1664 ();
 FILLCELL_X32 FILLCELL_208_1696 ();
 FILLCELL_X32 FILLCELL_208_1728 ();
 FILLCELL_X32 FILLCELL_208_1760 ();
 FILLCELL_X32 FILLCELL_208_1792 ();
 FILLCELL_X32 FILLCELL_208_1824 ();
 FILLCELL_X32 FILLCELL_208_1856 ();
 FILLCELL_X8 FILLCELL_208_1888 ();
 FILLCELL_X1 FILLCELL_208_1896 ();
 FILLCELL_X32 FILLCELL_209_0 ();
 FILLCELL_X32 FILLCELL_209_32 ();
 FILLCELL_X32 FILLCELL_209_64 ();
 FILLCELL_X32 FILLCELL_209_96 ();
 FILLCELL_X32 FILLCELL_209_128 ();
 FILLCELL_X32 FILLCELL_209_160 ();
 FILLCELL_X32 FILLCELL_209_192 ();
 FILLCELL_X32 FILLCELL_209_224 ();
 FILLCELL_X32 FILLCELL_209_256 ();
 FILLCELL_X32 FILLCELL_209_288 ();
 FILLCELL_X32 FILLCELL_209_320 ();
 FILLCELL_X32 FILLCELL_209_352 ();
 FILLCELL_X32 FILLCELL_209_384 ();
 FILLCELL_X32 FILLCELL_209_416 ();
 FILLCELL_X32 FILLCELL_209_448 ();
 FILLCELL_X32 FILLCELL_209_480 ();
 FILLCELL_X32 FILLCELL_209_512 ();
 FILLCELL_X32 FILLCELL_209_544 ();
 FILLCELL_X32 FILLCELL_209_576 ();
 FILLCELL_X32 FILLCELL_209_608 ();
 FILLCELL_X32 FILLCELL_209_640 ();
 FILLCELL_X32 FILLCELL_209_672 ();
 FILLCELL_X32 FILLCELL_209_704 ();
 FILLCELL_X32 FILLCELL_209_736 ();
 FILLCELL_X32 FILLCELL_209_768 ();
 FILLCELL_X32 FILLCELL_209_800 ();
 FILLCELL_X32 FILLCELL_209_832 ();
 FILLCELL_X32 FILLCELL_209_864 ();
 FILLCELL_X32 FILLCELL_209_896 ();
 FILLCELL_X32 FILLCELL_209_928 ();
 FILLCELL_X32 FILLCELL_209_960 ();
 FILLCELL_X32 FILLCELL_209_992 ();
 FILLCELL_X32 FILLCELL_209_1024 ();
 FILLCELL_X32 FILLCELL_209_1056 ();
 FILLCELL_X32 FILLCELL_209_1088 ();
 FILLCELL_X32 FILLCELL_209_1120 ();
 FILLCELL_X32 FILLCELL_209_1152 ();
 FILLCELL_X32 FILLCELL_209_1184 ();
 FILLCELL_X32 FILLCELL_209_1216 ();
 FILLCELL_X32 FILLCELL_209_1248 ();
 FILLCELL_X32 FILLCELL_209_1280 ();
 FILLCELL_X32 FILLCELL_209_1312 ();
 FILLCELL_X32 FILLCELL_209_1344 ();
 FILLCELL_X32 FILLCELL_209_1376 ();
 FILLCELL_X32 FILLCELL_209_1408 ();
 FILLCELL_X32 FILLCELL_209_1440 ();
 FILLCELL_X32 FILLCELL_209_1472 ();
 FILLCELL_X32 FILLCELL_209_1504 ();
 FILLCELL_X32 FILLCELL_209_1536 ();
 FILLCELL_X32 FILLCELL_209_1568 ();
 FILLCELL_X32 FILLCELL_209_1600 ();
 FILLCELL_X32 FILLCELL_209_1632 ();
 FILLCELL_X32 FILLCELL_209_1664 ();
 FILLCELL_X32 FILLCELL_209_1696 ();
 FILLCELL_X32 FILLCELL_209_1728 ();
 FILLCELL_X32 FILLCELL_209_1760 ();
 FILLCELL_X32 FILLCELL_209_1792 ();
 FILLCELL_X32 FILLCELL_209_1824 ();
 FILLCELL_X32 FILLCELL_209_1856 ();
 FILLCELL_X8 FILLCELL_209_1888 ();
 FILLCELL_X1 FILLCELL_209_1896 ();
 FILLCELL_X32 FILLCELL_210_0 ();
 FILLCELL_X32 FILLCELL_210_32 ();
 FILLCELL_X32 FILLCELL_210_64 ();
 FILLCELL_X32 FILLCELL_210_96 ();
 FILLCELL_X32 FILLCELL_210_128 ();
 FILLCELL_X32 FILLCELL_210_160 ();
 FILLCELL_X32 FILLCELL_210_192 ();
 FILLCELL_X32 FILLCELL_210_224 ();
 FILLCELL_X32 FILLCELL_210_256 ();
 FILLCELL_X32 FILLCELL_210_288 ();
 FILLCELL_X32 FILLCELL_210_320 ();
 FILLCELL_X32 FILLCELL_210_352 ();
 FILLCELL_X32 FILLCELL_210_384 ();
 FILLCELL_X32 FILLCELL_210_416 ();
 FILLCELL_X32 FILLCELL_210_448 ();
 FILLCELL_X32 FILLCELL_210_480 ();
 FILLCELL_X32 FILLCELL_210_512 ();
 FILLCELL_X32 FILLCELL_210_544 ();
 FILLCELL_X32 FILLCELL_210_576 ();
 FILLCELL_X32 FILLCELL_210_608 ();
 FILLCELL_X32 FILLCELL_210_640 ();
 FILLCELL_X32 FILLCELL_210_672 ();
 FILLCELL_X32 FILLCELL_210_704 ();
 FILLCELL_X32 FILLCELL_210_736 ();
 FILLCELL_X32 FILLCELL_210_768 ();
 FILLCELL_X32 FILLCELL_210_800 ();
 FILLCELL_X32 FILLCELL_210_832 ();
 FILLCELL_X32 FILLCELL_210_864 ();
 FILLCELL_X32 FILLCELL_210_896 ();
 FILLCELL_X32 FILLCELL_210_928 ();
 FILLCELL_X32 FILLCELL_210_960 ();
 FILLCELL_X32 FILLCELL_210_992 ();
 FILLCELL_X32 FILLCELL_210_1024 ();
 FILLCELL_X32 FILLCELL_210_1056 ();
 FILLCELL_X32 FILLCELL_210_1088 ();
 FILLCELL_X32 FILLCELL_210_1120 ();
 FILLCELL_X32 FILLCELL_210_1152 ();
 FILLCELL_X32 FILLCELL_210_1184 ();
 FILLCELL_X32 FILLCELL_210_1216 ();
 FILLCELL_X32 FILLCELL_210_1248 ();
 FILLCELL_X32 FILLCELL_210_1280 ();
 FILLCELL_X32 FILLCELL_210_1312 ();
 FILLCELL_X32 FILLCELL_210_1344 ();
 FILLCELL_X32 FILLCELL_210_1376 ();
 FILLCELL_X32 FILLCELL_210_1408 ();
 FILLCELL_X32 FILLCELL_210_1440 ();
 FILLCELL_X32 FILLCELL_210_1472 ();
 FILLCELL_X32 FILLCELL_210_1504 ();
 FILLCELL_X32 FILLCELL_210_1536 ();
 FILLCELL_X32 FILLCELL_210_1568 ();
 FILLCELL_X32 FILLCELL_210_1600 ();
 FILLCELL_X32 FILLCELL_210_1632 ();
 FILLCELL_X32 FILLCELL_210_1664 ();
 FILLCELL_X32 FILLCELL_210_1696 ();
 FILLCELL_X32 FILLCELL_210_1728 ();
 FILLCELL_X32 FILLCELL_210_1760 ();
 FILLCELL_X32 FILLCELL_210_1792 ();
 FILLCELL_X32 FILLCELL_210_1824 ();
 FILLCELL_X32 FILLCELL_210_1856 ();
 FILLCELL_X8 FILLCELL_210_1888 ();
 FILLCELL_X1 FILLCELL_210_1896 ();
 FILLCELL_X32 FILLCELL_211_0 ();
 FILLCELL_X32 FILLCELL_211_32 ();
 FILLCELL_X32 FILLCELL_211_64 ();
 FILLCELL_X32 FILLCELL_211_96 ();
 FILLCELL_X32 FILLCELL_211_128 ();
 FILLCELL_X32 FILLCELL_211_160 ();
 FILLCELL_X32 FILLCELL_211_192 ();
 FILLCELL_X32 FILLCELL_211_224 ();
 FILLCELL_X32 FILLCELL_211_256 ();
 FILLCELL_X32 FILLCELL_211_288 ();
 FILLCELL_X32 FILLCELL_211_320 ();
 FILLCELL_X32 FILLCELL_211_352 ();
 FILLCELL_X32 FILLCELL_211_384 ();
 FILLCELL_X32 FILLCELL_211_416 ();
 FILLCELL_X32 FILLCELL_211_448 ();
 FILLCELL_X32 FILLCELL_211_480 ();
 FILLCELL_X32 FILLCELL_211_512 ();
 FILLCELL_X32 FILLCELL_211_544 ();
 FILLCELL_X32 FILLCELL_211_576 ();
 FILLCELL_X32 FILLCELL_211_608 ();
 FILLCELL_X32 FILLCELL_211_640 ();
 FILLCELL_X32 FILLCELL_211_672 ();
 FILLCELL_X32 FILLCELL_211_704 ();
 FILLCELL_X32 FILLCELL_211_736 ();
 FILLCELL_X32 FILLCELL_211_768 ();
 FILLCELL_X32 FILLCELL_211_800 ();
 FILLCELL_X32 FILLCELL_211_832 ();
 FILLCELL_X32 FILLCELL_211_864 ();
 FILLCELL_X32 FILLCELL_211_896 ();
 FILLCELL_X32 FILLCELL_211_928 ();
 FILLCELL_X32 FILLCELL_211_960 ();
 FILLCELL_X32 FILLCELL_211_992 ();
 FILLCELL_X32 FILLCELL_211_1024 ();
 FILLCELL_X32 FILLCELL_211_1056 ();
 FILLCELL_X32 FILLCELL_211_1088 ();
 FILLCELL_X32 FILLCELL_211_1120 ();
 FILLCELL_X32 FILLCELL_211_1152 ();
 FILLCELL_X32 FILLCELL_211_1184 ();
 FILLCELL_X32 FILLCELL_211_1216 ();
 FILLCELL_X32 FILLCELL_211_1248 ();
 FILLCELL_X32 FILLCELL_211_1280 ();
 FILLCELL_X32 FILLCELL_211_1312 ();
 FILLCELL_X32 FILLCELL_211_1344 ();
 FILLCELL_X32 FILLCELL_211_1376 ();
 FILLCELL_X32 FILLCELL_211_1408 ();
 FILLCELL_X32 FILLCELL_211_1440 ();
 FILLCELL_X32 FILLCELL_211_1472 ();
 FILLCELL_X32 FILLCELL_211_1504 ();
 FILLCELL_X32 FILLCELL_211_1536 ();
 FILLCELL_X32 FILLCELL_211_1568 ();
 FILLCELL_X32 FILLCELL_211_1600 ();
 FILLCELL_X32 FILLCELL_211_1632 ();
 FILLCELL_X32 FILLCELL_211_1664 ();
 FILLCELL_X32 FILLCELL_211_1696 ();
 FILLCELL_X32 FILLCELL_211_1728 ();
 FILLCELL_X32 FILLCELL_211_1760 ();
 FILLCELL_X32 FILLCELL_211_1792 ();
 FILLCELL_X32 FILLCELL_211_1824 ();
 FILLCELL_X32 FILLCELL_211_1856 ();
 FILLCELL_X8 FILLCELL_211_1888 ();
 FILLCELL_X1 FILLCELL_211_1896 ();
 FILLCELL_X32 FILLCELL_212_0 ();
 FILLCELL_X32 FILLCELL_212_32 ();
 FILLCELL_X32 FILLCELL_212_64 ();
 FILLCELL_X32 FILLCELL_212_96 ();
 FILLCELL_X32 FILLCELL_212_128 ();
 FILLCELL_X32 FILLCELL_212_160 ();
 FILLCELL_X32 FILLCELL_212_192 ();
 FILLCELL_X32 FILLCELL_212_224 ();
 FILLCELL_X32 FILLCELL_212_256 ();
 FILLCELL_X32 FILLCELL_212_288 ();
 FILLCELL_X32 FILLCELL_212_320 ();
 FILLCELL_X32 FILLCELL_212_352 ();
 FILLCELL_X32 FILLCELL_212_384 ();
 FILLCELL_X32 FILLCELL_212_416 ();
 FILLCELL_X32 FILLCELL_212_448 ();
 FILLCELL_X32 FILLCELL_212_480 ();
 FILLCELL_X32 FILLCELL_212_512 ();
 FILLCELL_X32 FILLCELL_212_544 ();
 FILLCELL_X32 FILLCELL_212_576 ();
 FILLCELL_X32 FILLCELL_212_608 ();
 FILLCELL_X32 FILLCELL_212_640 ();
 FILLCELL_X32 FILLCELL_212_672 ();
 FILLCELL_X32 FILLCELL_212_704 ();
 FILLCELL_X32 FILLCELL_212_736 ();
 FILLCELL_X32 FILLCELL_212_768 ();
 FILLCELL_X32 FILLCELL_212_800 ();
 FILLCELL_X32 FILLCELL_212_832 ();
 FILLCELL_X32 FILLCELL_212_864 ();
 FILLCELL_X32 FILLCELL_212_896 ();
 FILLCELL_X32 FILLCELL_212_928 ();
 FILLCELL_X32 FILLCELL_212_960 ();
 FILLCELL_X32 FILLCELL_212_992 ();
 FILLCELL_X32 FILLCELL_212_1024 ();
 FILLCELL_X32 FILLCELL_212_1056 ();
 FILLCELL_X32 FILLCELL_212_1088 ();
 FILLCELL_X32 FILLCELL_212_1120 ();
 FILLCELL_X32 FILLCELL_212_1152 ();
 FILLCELL_X32 FILLCELL_212_1184 ();
 FILLCELL_X32 FILLCELL_212_1216 ();
 FILLCELL_X32 FILLCELL_212_1248 ();
 FILLCELL_X32 FILLCELL_212_1280 ();
 FILLCELL_X32 FILLCELL_212_1312 ();
 FILLCELL_X32 FILLCELL_212_1344 ();
 FILLCELL_X32 FILLCELL_212_1376 ();
 FILLCELL_X32 FILLCELL_212_1408 ();
 FILLCELL_X32 FILLCELL_212_1440 ();
 FILLCELL_X32 FILLCELL_212_1472 ();
 FILLCELL_X32 FILLCELL_212_1504 ();
 FILLCELL_X32 FILLCELL_212_1536 ();
 FILLCELL_X32 FILLCELL_212_1568 ();
 FILLCELL_X32 FILLCELL_212_1600 ();
 FILLCELL_X32 FILLCELL_212_1632 ();
 FILLCELL_X32 FILLCELL_212_1664 ();
 FILLCELL_X32 FILLCELL_212_1696 ();
 FILLCELL_X32 FILLCELL_212_1728 ();
 FILLCELL_X32 FILLCELL_212_1760 ();
 FILLCELL_X32 FILLCELL_212_1792 ();
 FILLCELL_X32 FILLCELL_212_1824 ();
 FILLCELL_X32 FILLCELL_212_1856 ();
 FILLCELL_X8 FILLCELL_212_1888 ();
 FILLCELL_X1 FILLCELL_212_1896 ();
 FILLCELL_X32 FILLCELL_213_0 ();
 FILLCELL_X32 FILLCELL_213_32 ();
 FILLCELL_X32 FILLCELL_213_64 ();
 FILLCELL_X32 FILLCELL_213_96 ();
 FILLCELL_X32 FILLCELL_213_128 ();
 FILLCELL_X32 FILLCELL_213_160 ();
 FILLCELL_X32 FILLCELL_213_192 ();
 FILLCELL_X32 FILLCELL_213_224 ();
 FILLCELL_X32 FILLCELL_213_256 ();
 FILLCELL_X32 FILLCELL_213_288 ();
 FILLCELL_X32 FILLCELL_213_320 ();
 FILLCELL_X32 FILLCELL_213_352 ();
 FILLCELL_X32 FILLCELL_213_384 ();
 FILLCELL_X32 FILLCELL_213_416 ();
 FILLCELL_X32 FILLCELL_213_448 ();
 FILLCELL_X32 FILLCELL_213_480 ();
 FILLCELL_X32 FILLCELL_213_512 ();
 FILLCELL_X32 FILLCELL_213_544 ();
 FILLCELL_X32 FILLCELL_213_576 ();
 FILLCELL_X32 FILLCELL_213_608 ();
 FILLCELL_X32 FILLCELL_213_640 ();
 FILLCELL_X32 FILLCELL_213_672 ();
 FILLCELL_X32 FILLCELL_213_704 ();
 FILLCELL_X32 FILLCELL_213_736 ();
 FILLCELL_X32 FILLCELL_213_768 ();
 FILLCELL_X32 FILLCELL_213_800 ();
 FILLCELL_X32 FILLCELL_213_832 ();
 FILLCELL_X32 FILLCELL_213_864 ();
 FILLCELL_X32 FILLCELL_213_896 ();
 FILLCELL_X32 FILLCELL_213_928 ();
 FILLCELL_X32 FILLCELL_213_960 ();
 FILLCELL_X32 FILLCELL_213_992 ();
 FILLCELL_X32 FILLCELL_213_1024 ();
 FILLCELL_X32 FILLCELL_213_1056 ();
 FILLCELL_X32 FILLCELL_213_1088 ();
 FILLCELL_X32 FILLCELL_213_1120 ();
 FILLCELL_X32 FILLCELL_213_1152 ();
 FILLCELL_X32 FILLCELL_213_1184 ();
 FILLCELL_X32 FILLCELL_213_1216 ();
 FILLCELL_X32 FILLCELL_213_1248 ();
 FILLCELL_X32 FILLCELL_213_1280 ();
 FILLCELL_X32 FILLCELL_213_1312 ();
 FILLCELL_X32 FILLCELL_213_1344 ();
 FILLCELL_X32 FILLCELL_213_1376 ();
 FILLCELL_X32 FILLCELL_213_1408 ();
 FILLCELL_X32 FILLCELL_213_1440 ();
 FILLCELL_X32 FILLCELL_213_1472 ();
 FILLCELL_X32 FILLCELL_213_1504 ();
 FILLCELL_X32 FILLCELL_213_1536 ();
 FILLCELL_X32 FILLCELL_213_1568 ();
 FILLCELL_X32 FILLCELL_213_1600 ();
 FILLCELL_X32 FILLCELL_213_1632 ();
 FILLCELL_X32 FILLCELL_213_1664 ();
 FILLCELL_X32 FILLCELL_213_1696 ();
 FILLCELL_X32 FILLCELL_213_1728 ();
 FILLCELL_X32 FILLCELL_213_1760 ();
 FILLCELL_X32 FILLCELL_213_1792 ();
 FILLCELL_X32 FILLCELL_213_1824 ();
 FILLCELL_X32 FILLCELL_213_1856 ();
 FILLCELL_X8 FILLCELL_213_1888 ();
 FILLCELL_X1 FILLCELL_213_1896 ();
 FILLCELL_X32 FILLCELL_214_0 ();
 FILLCELL_X32 FILLCELL_214_32 ();
 FILLCELL_X32 FILLCELL_214_64 ();
 FILLCELL_X32 FILLCELL_214_96 ();
 FILLCELL_X32 FILLCELL_214_128 ();
 FILLCELL_X32 FILLCELL_214_160 ();
 FILLCELL_X32 FILLCELL_214_192 ();
 FILLCELL_X32 FILLCELL_214_224 ();
 FILLCELL_X32 FILLCELL_214_256 ();
 FILLCELL_X32 FILLCELL_214_288 ();
 FILLCELL_X32 FILLCELL_214_320 ();
 FILLCELL_X32 FILLCELL_214_352 ();
 FILLCELL_X32 FILLCELL_214_384 ();
 FILLCELL_X32 FILLCELL_214_416 ();
 FILLCELL_X32 FILLCELL_214_448 ();
 FILLCELL_X32 FILLCELL_214_480 ();
 FILLCELL_X32 FILLCELL_214_512 ();
 FILLCELL_X32 FILLCELL_214_544 ();
 FILLCELL_X32 FILLCELL_214_576 ();
 FILLCELL_X32 FILLCELL_214_608 ();
 FILLCELL_X32 FILLCELL_214_640 ();
 FILLCELL_X32 FILLCELL_214_672 ();
 FILLCELL_X32 FILLCELL_214_704 ();
 FILLCELL_X32 FILLCELL_214_736 ();
 FILLCELL_X32 FILLCELL_214_768 ();
 FILLCELL_X32 FILLCELL_214_800 ();
 FILLCELL_X32 FILLCELL_214_832 ();
 FILLCELL_X32 FILLCELL_214_864 ();
 FILLCELL_X32 FILLCELL_214_896 ();
 FILLCELL_X32 FILLCELL_214_928 ();
 FILLCELL_X32 FILLCELL_214_960 ();
 FILLCELL_X32 FILLCELL_214_992 ();
 FILLCELL_X32 FILLCELL_214_1024 ();
 FILLCELL_X32 FILLCELL_214_1056 ();
 FILLCELL_X32 FILLCELL_214_1088 ();
 FILLCELL_X32 FILLCELL_214_1120 ();
 FILLCELL_X32 FILLCELL_214_1152 ();
 FILLCELL_X32 FILLCELL_214_1184 ();
 FILLCELL_X32 FILLCELL_214_1216 ();
 FILLCELL_X32 FILLCELL_214_1248 ();
 FILLCELL_X32 FILLCELL_214_1280 ();
 FILLCELL_X32 FILLCELL_214_1312 ();
 FILLCELL_X32 FILLCELL_214_1344 ();
 FILLCELL_X32 FILLCELL_214_1376 ();
 FILLCELL_X32 FILLCELL_214_1408 ();
 FILLCELL_X32 FILLCELL_214_1440 ();
 FILLCELL_X32 FILLCELL_214_1472 ();
 FILLCELL_X32 FILLCELL_214_1504 ();
 FILLCELL_X32 FILLCELL_214_1536 ();
 FILLCELL_X32 FILLCELL_214_1568 ();
 FILLCELL_X32 FILLCELL_214_1600 ();
 FILLCELL_X32 FILLCELL_214_1632 ();
 FILLCELL_X32 FILLCELL_214_1664 ();
 FILLCELL_X32 FILLCELL_214_1696 ();
 FILLCELL_X32 FILLCELL_214_1728 ();
 FILLCELL_X32 FILLCELL_214_1760 ();
 FILLCELL_X32 FILLCELL_214_1792 ();
 FILLCELL_X32 FILLCELL_214_1824 ();
 FILLCELL_X32 FILLCELL_214_1856 ();
 FILLCELL_X8 FILLCELL_214_1888 ();
 FILLCELL_X1 FILLCELL_214_1896 ();
 FILLCELL_X32 FILLCELL_215_0 ();
 FILLCELL_X32 FILLCELL_215_32 ();
 FILLCELL_X32 FILLCELL_215_64 ();
 FILLCELL_X32 FILLCELL_215_96 ();
 FILLCELL_X32 FILLCELL_215_128 ();
 FILLCELL_X32 FILLCELL_215_160 ();
 FILLCELL_X32 FILLCELL_215_192 ();
 FILLCELL_X32 FILLCELL_215_224 ();
 FILLCELL_X32 FILLCELL_215_256 ();
 FILLCELL_X32 FILLCELL_215_288 ();
 FILLCELL_X32 FILLCELL_215_320 ();
 FILLCELL_X32 FILLCELL_215_352 ();
 FILLCELL_X32 FILLCELL_215_384 ();
 FILLCELL_X32 FILLCELL_215_416 ();
 FILLCELL_X32 FILLCELL_215_448 ();
 FILLCELL_X32 FILLCELL_215_480 ();
 FILLCELL_X32 FILLCELL_215_512 ();
 FILLCELL_X32 FILLCELL_215_544 ();
 FILLCELL_X32 FILLCELL_215_576 ();
 FILLCELL_X32 FILLCELL_215_608 ();
 FILLCELL_X32 FILLCELL_215_640 ();
 FILLCELL_X32 FILLCELL_215_672 ();
 FILLCELL_X32 FILLCELL_215_704 ();
 FILLCELL_X32 FILLCELL_215_736 ();
 FILLCELL_X32 FILLCELL_215_768 ();
 FILLCELL_X32 FILLCELL_215_800 ();
 FILLCELL_X32 FILLCELL_215_832 ();
 FILLCELL_X32 FILLCELL_215_864 ();
 FILLCELL_X32 FILLCELL_215_896 ();
 FILLCELL_X32 FILLCELL_215_928 ();
 FILLCELL_X32 FILLCELL_215_960 ();
 FILLCELL_X32 FILLCELL_215_992 ();
 FILLCELL_X32 FILLCELL_215_1024 ();
 FILLCELL_X32 FILLCELL_215_1056 ();
 FILLCELL_X32 FILLCELL_215_1088 ();
 FILLCELL_X32 FILLCELL_215_1120 ();
 FILLCELL_X32 FILLCELL_215_1152 ();
 FILLCELL_X32 FILLCELL_215_1184 ();
 FILLCELL_X32 FILLCELL_215_1216 ();
 FILLCELL_X32 FILLCELL_215_1248 ();
 FILLCELL_X32 FILLCELL_215_1280 ();
 FILLCELL_X32 FILLCELL_215_1312 ();
 FILLCELL_X32 FILLCELL_215_1344 ();
 FILLCELL_X32 FILLCELL_215_1376 ();
 FILLCELL_X32 FILLCELL_215_1408 ();
 FILLCELL_X32 FILLCELL_215_1440 ();
 FILLCELL_X32 FILLCELL_215_1472 ();
 FILLCELL_X32 FILLCELL_215_1504 ();
 FILLCELL_X32 FILLCELL_215_1536 ();
 FILLCELL_X32 FILLCELL_215_1568 ();
 FILLCELL_X32 FILLCELL_215_1600 ();
 FILLCELL_X32 FILLCELL_215_1632 ();
 FILLCELL_X32 FILLCELL_215_1664 ();
 FILLCELL_X32 FILLCELL_215_1696 ();
 FILLCELL_X32 FILLCELL_215_1728 ();
 FILLCELL_X32 FILLCELL_215_1760 ();
 FILLCELL_X32 FILLCELL_215_1792 ();
 FILLCELL_X32 FILLCELL_215_1824 ();
 FILLCELL_X32 FILLCELL_215_1856 ();
 FILLCELL_X8 FILLCELL_215_1888 ();
 FILLCELL_X1 FILLCELL_215_1896 ();
 FILLCELL_X32 FILLCELL_216_0 ();
 FILLCELL_X32 FILLCELL_216_32 ();
 FILLCELL_X32 FILLCELL_216_64 ();
 FILLCELL_X32 FILLCELL_216_96 ();
 FILLCELL_X32 FILLCELL_216_128 ();
 FILLCELL_X32 FILLCELL_216_160 ();
 FILLCELL_X32 FILLCELL_216_192 ();
 FILLCELL_X32 FILLCELL_216_224 ();
 FILLCELL_X32 FILLCELL_216_256 ();
 FILLCELL_X32 FILLCELL_216_288 ();
 FILLCELL_X32 FILLCELL_216_320 ();
 FILLCELL_X32 FILLCELL_216_352 ();
 FILLCELL_X32 FILLCELL_216_384 ();
 FILLCELL_X32 FILLCELL_216_416 ();
 FILLCELL_X32 FILLCELL_216_448 ();
 FILLCELL_X32 FILLCELL_216_480 ();
 FILLCELL_X32 FILLCELL_216_512 ();
 FILLCELL_X32 FILLCELL_216_544 ();
 FILLCELL_X32 FILLCELL_216_576 ();
 FILLCELL_X32 FILLCELL_216_608 ();
 FILLCELL_X32 FILLCELL_216_640 ();
 FILLCELL_X32 FILLCELL_216_672 ();
 FILLCELL_X32 FILLCELL_216_704 ();
 FILLCELL_X32 FILLCELL_216_736 ();
 FILLCELL_X32 FILLCELL_216_768 ();
 FILLCELL_X32 FILLCELL_216_800 ();
 FILLCELL_X32 FILLCELL_216_832 ();
 FILLCELL_X32 FILLCELL_216_864 ();
 FILLCELL_X32 FILLCELL_216_896 ();
 FILLCELL_X32 FILLCELL_216_928 ();
 FILLCELL_X32 FILLCELL_216_960 ();
 FILLCELL_X32 FILLCELL_216_992 ();
 FILLCELL_X32 FILLCELL_216_1024 ();
 FILLCELL_X32 FILLCELL_216_1056 ();
 FILLCELL_X32 FILLCELL_216_1088 ();
 FILLCELL_X32 FILLCELL_216_1120 ();
 FILLCELL_X32 FILLCELL_216_1152 ();
 FILLCELL_X32 FILLCELL_216_1184 ();
 FILLCELL_X32 FILLCELL_216_1216 ();
 FILLCELL_X32 FILLCELL_216_1248 ();
 FILLCELL_X32 FILLCELL_216_1280 ();
 FILLCELL_X32 FILLCELL_216_1312 ();
 FILLCELL_X32 FILLCELL_216_1344 ();
 FILLCELL_X32 FILLCELL_216_1376 ();
 FILLCELL_X32 FILLCELL_216_1408 ();
 FILLCELL_X32 FILLCELL_216_1440 ();
 FILLCELL_X32 FILLCELL_216_1472 ();
 FILLCELL_X32 FILLCELL_216_1504 ();
 FILLCELL_X32 FILLCELL_216_1536 ();
 FILLCELL_X32 FILLCELL_216_1568 ();
 FILLCELL_X32 FILLCELL_216_1600 ();
 FILLCELL_X32 FILLCELL_216_1632 ();
 FILLCELL_X32 FILLCELL_216_1664 ();
 FILLCELL_X32 FILLCELL_216_1696 ();
 FILLCELL_X32 FILLCELL_216_1728 ();
 FILLCELL_X32 FILLCELL_216_1760 ();
 FILLCELL_X32 FILLCELL_216_1792 ();
 FILLCELL_X32 FILLCELL_216_1824 ();
 FILLCELL_X32 FILLCELL_216_1856 ();
 FILLCELL_X8 FILLCELL_216_1888 ();
 FILLCELL_X1 FILLCELL_216_1896 ();
 FILLCELL_X32 FILLCELL_217_0 ();
 FILLCELL_X32 FILLCELL_217_32 ();
 FILLCELL_X32 FILLCELL_217_64 ();
 FILLCELL_X32 FILLCELL_217_96 ();
 FILLCELL_X32 FILLCELL_217_128 ();
 FILLCELL_X32 FILLCELL_217_160 ();
 FILLCELL_X32 FILLCELL_217_192 ();
 FILLCELL_X32 FILLCELL_217_224 ();
 FILLCELL_X32 FILLCELL_217_256 ();
 FILLCELL_X32 FILLCELL_217_288 ();
 FILLCELL_X32 FILLCELL_217_320 ();
 FILLCELL_X32 FILLCELL_217_352 ();
 FILLCELL_X32 FILLCELL_217_384 ();
 FILLCELL_X32 FILLCELL_217_416 ();
 FILLCELL_X32 FILLCELL_217_448 ();
 FILLCELL_X32 FILLCELL_217_480 ();
 FILLCELL_X32 FILLCELL_217_512 ();
 FILLCELL_X32 FILLCELL_217_544 ();
 FILLCELL_X32 FILLCELL_217_576 ();
 FILLCELL_X32 FILLCELL_217_608 ();
 FILLCELL_X32 FILLCELL_217_640 ();
 FILLCELL_X32 FILLCELL_217_672 ();
 FILLCELL_X32 FILLCELL_217_704 ();
 FILLCELL_X32 FILLCELL_217_736 ();
 FILLCELL_X32 FILLCELL_217_768 ();
 FILLCELL_X32 FILLCELL_217_800 ();
 FILLCELL_X32 FILLCELL_217_832 ();
 FILLCELL_X32 FILLCELL_217_864 ();
 FILLCELL_X32 FILLCELL_217_896 ();
 FILLCELL_X32 FILLCELL_217_928 ();
 FILLCELL_X32 FILLCELL_217_960 ();
 FILLCELL_X32 FILLCELL_217_992 ();
 FILLCELL_X32 FILLCELL_217_1024 ();
 FILLCELL_X32 FILLCELL_217_1056 ();
 FILLCELL_X32 FILLCELL_217_1088 ();
 FILLCELL_X32 FILLCELL_217_1120 ();
 FILLCELL_X32 FILLCELL_217_1152 ();
 FILLCELL_X32 FILLCELL_217_1184 ();
 FILLCELL_X32 FILLCELL_217_1216 ();
 FILLCELL_X32 FILLCELL_217_1248 ();
 FILLCELL_X32 FILLCELL_217_1280 ();
 FILLCELL_X32 FILLCELL_217_1312 ();
 FILLCELL_X32 FILLCELL_217_1344 ();
 FILLCELL_X32 FILLCELL_217_1376 ();
 FILLCELL_X32 FILLCELL_217_1408 ();
 FILLCELL_X32 FILLCELL_217_1440 ();
 FILLCELL_X32 FILLCELL_217_1472 ();
 FILLCELL_X32 FILLCELL_217_1504 ();
 FILLCELL_X32 FILLCELL_217_1536 ();
 FILLCELL_X32 FILLCELL_217_1568 ();
 FILLCELL_X32 FILLCELL_217_1600 ();
 FILLCELL_X32 FILLCELL_217_1632 ();
 FILLCELL_X32 FILLCELL_217_1664 ();
 FILLCELL_X32 FILLCELL_217_1696 ();
 FILLCELL_X32 FILLCELL_217_1728 ();
 FILLCELL_X32 FILLCELL_217_1760 ();
 FILLCELL_X32 FILLCELL_217_1792 ();
 FILLCELL_X32 FILLCELL_217_1824 ();
 FILLCELL_X32 FILLCELL_217_1856 ();
 FILLCELL_X8 FILLCELL_217_1888 ();
 FILLCELL_X1 FILLCELL_217_1896 ();
 FILLCELL_X32 FILLCELL_218_0 ();
 FILLCELL_X32 FILLCELL_218_32 ();
 FILLCELL_X32 FILLCELL_218_64 ();
 FILLCELL_X32 FILLCELL_218_96 ();
 FILLCELL_X32 FILLCELL_218_128 ();
 FILLCELL_X32 FILLCELL_218_160 ();
 FILLCELL_X32 FILLCELL_218_192 ();
 FILLCELL_X32 FILLCELL_218_224 ();
 FILLCELL_X32 FILLCELL_218_256 ();
 FILLCELL_X32 FILLCELL_218_288 ();
 FILLCELL_X32 FILLCELL_218_320 ();
 FILLCELL_X32 FILLCELL_218_352 ();
 FILLCELL_X32 FILLCELL_218_384 ();
 FILLCELL_X32 FILLCELL_218_416 ();
 FILLCELL_X32 FILLCELL_218_448 ();
 FILLCELL_X32 FILLCELL_218_480 ();
 FILLCELL_X32 FILLCELL_218_512 ();
 FILLCELL_X32 FILLCELL_218_544 ();
 FILLCELL_X32 FILLCELL_218_576 ();
 FILLCELL_X32 FILLCELL_218_608 ();
 FILLCELL_X32 FILLCELL_218_640 ();
 FILLCELL_X32 FILLCELL_218_672 ();
 FILLCELL_X32 FILLCELL_218_704 ();
 FILLCELL_X32 FILLCELL_218_736 ();
 FILLCELL_X32 FILLCELL_218_768 ();
 FILLCELL_X32 FILLCELL_218_800 ();
 FILLCELL_X32 FILLCELL_218_832 ();
 FILLCELL_X32 FILLCELL_218_864 ();
 FILLCELL_X32 FILLCELL_218_896 ();
 FILLCELL_X32 FILLCELL_218_928 ();
 FILLCELL_X32 FILLCELL_218_960 ();
 FILLCELL_X32 FILLCELL_218_992 ();
 FILLCELL_X32 FILLCELL_218_1024 ();
 FILLCELL_X32 FILLCELL_218_1056 ();
 FILLCELL_X32 FILLCELL_218_1088 ();
 FILLCELL_X32 FILLCELL_218_1120 ();
 FILLCELL_X32 FILLCELL_218_1152 ();
 FILLCELL_X32 FILLCELL_218_1184 ();
 FILLCELL_X32 FILLCELL_218_1216 ();
 FILLCELL_X32 FILLCELL_218_1248 ();
 FILLCELL_X32 FILLCELL_218_1280 ();
 FILLCELL_X32 FILLCELL_218_1312 ();
 FILLCELL_X32 FILLCELL_218_1344 ();
 FILLCELL_X32 FILLCELL_218_1376 ();
 FILLCELL_X32 FILLCELL_218_1408 ();
 FILLCELL_X32 FILLCELL_218_1440 ();
 FILLCELL_X32 FILLCELL_218_1472 ();
 FILLCELL_X32 FILLCELL_218_1504 ();
 FILLCELL_X32 FILLCELL_218_1536 ();
 FILLCELL_X32 FILLCELL_218_1568 ();
 FILLCELL_X32 FILLCELL_218_1600 ();
 FILLCELL_X32 FILLCELL_218_1632 ();
 FILLCELL_X32 FILLCELL_218_1664 ();
 FILLCELL_X32 FILLCELL_218_1696 ();
 FILLCELL_X32 FILLCELL_218_1728 ();
 FILLCELL_X32 FILLCELL_218_1760 ();
 FILLCELL_X32 FILLCELL_218_1792 ();
 FILLCELL_X32 FILLCELL_218_1824 ();
 FILLCELL_X32 FILLCELL_218_1856 ();
 FILLCELL_X8 FILLCELL_218_1888 ();
 FILLCELL_X1 FILLCELL_218_1896 ();
 FILLCELL_X32 FILLCELL_219_0 ();
 FILLCELL_X32 FILLCELL_219_32 ();
 FILLCELL_X32 FILLCELL_219_64 ();
 FILLCELL_X32 FILLCELL_219_96 ();
 FILLCELL_X32 FILLCELL_219_128 ();
 FILLCELL_X32 FILLCELL_219_160 ();
 FILLCELL_X32 FILLCELL_219_192 ();
 FILLCELL_X32 FILLCELL_219_224 ();
 FILLCELL_X32 FILLCELL_219_256 ();
 FILLCELL_X32 FILLCELL_219_288 ();
 FILLCELL_X32 FILLCELL_219_320 ();
 FILLCELL_X32 FILLCELL_219_352 ();
 FILLCELL_X32 FILLCELL_219_384 ();
 FILLCELL_X32 FILLCELL_219_416 ();
 FILLCELL_X32 FILLCELL_219_448 ();
 FILLCELL_X32 FILLCELL_219_480 ();
 FILLCELL_X32 FILLCELL_219_512 ();
 FILLCELL_X32 FILLCELL_219_544 ();
 FILLCELL_X32 FILLCELL_219_576 ();
 FILLCELL_X32 FILLCELL_219_608 ();
 FILLCELL_X32 FILLCELL_219_640 ();
 FILLCELL_X32 FILLCELL_219_672 ();
 FILLCELL_X32 FILLCELL_219_704 ();
 FILLCELL_X32 FILLCELL_219_736 ();
 FILLCELL_X32 FILLCELL_219_768 ();
 FILLCELL_X32 FILLCELL_219_800 ();
 FILLCELL_X32 FILLCELL_219_832 ();
 FILLCELL_X32 FILLCELL_219_864 ();
 FILLCELL_X32 FILLCELL_219_896 ();
 FILLCELL_X32 FILLCELL_219_928 ();
 FILLCELL_X32 FILLCELL_219_960 ();
 FILLCELL_X32 FILLCELL_219_992 ();
 FILLCELL_X32 FILLCELL_219_1024 ();
 FILLCELL_X32 FILLCELL_219_1056 ();
 FILLCELL_X32 FILLCELL_219_1088 ();
 FILLCELL_X32 FILLCELL_219_1120 ();
 FILLCELL_X32 FILLCELL_219_1152 ();
 FILLCELL_X32 FILLCELL_219_1184 ();
 FILLCELL_X32 FILLCELL_219_1216 ();
 FILLCELL_X32 FILLCELL_219_1248 ();
 FILLCELL_X32 FILLCELL_219_1280 ();
 FILLCELL_X32 FILLCELL_219_1312 ();
 FILLCELL_X32 FILLCELL_219_1344 ();
 FILLCELL_X32 FILLCELL_219_1376 ();
 FILLCELL_X32 FILLCELL_219_1408 ();
 FILLCELL_X32 FILLCELL_219_1440 ();
 FILLCELL_X32 FILLCELL_219_1472 ();
 FILLCELL_X32 FILLCELL_219_1504 ();
 FILLCELL_X32 FILLCELL_219_1536 ();
 FILLCELL_X32 FILLCELL_219_1568 ();
 FILLCELL_X32 FILLCELL_219_1600 ();
 FILLCELL_X32 FILLCELL_219_1632 ();
 FILLCELL_X32 FILLCELL_219_1664 ();
 FILLCELL_X32 FILLCELL_219_1696 ();
 FILLCELL_X32 FILLCELL_219_1728 ();
 FILLCELL_X32 FILLCELL_219_1760 ();
 FILLCELL_X32 FILLCELL_219_1792 ();
 FILLCELL_X32 FILLCELL_219_1824 ();
 FILLCELL_X32 FILLCELL_219_1856 ();
 FILLCELL_X8 FILLCELL_219_1888 ();
 FILLCELL_X1 FILLCELL_219_1896 ();
 FILLCELL_X32 FILLCELL_220_0 ();
 FILLCELL_X32 FILLCELL_220_32 ();
 FILLCELL_X32 FILLCELL_220_64 ();
 FILLCELL_X32 FILLCELL_220_96 ();
 FILLCELL_X32 FILLCELL_220_128 ();
 FILLCELL_X32 FILLCELL_220_160 ();
 FILLCELL_X32 FILLCELL_220_192 ();
 FILLCELL_X32 FILLCELL_220_224 ();
 FILLCELL_X32 FILLCELL_220_256 ();
 FILLCELL_X32 FILLCELL_220_288 ();
 FILLCELL_X32 FILLCELL_220_320 ();
 FILLCELL_X32 FILLCELL_220_352 ();
 FILLCELL_X32 FILLCELL_220_384 ();
 FILLCELL_X32 FILLCELL_220_416 ();
 FILLCELL_X32 FILLCELL_220_448 ();
 FILLCELL_X32 FILLCELL_220_480 ();
 FILLCELL_X32 FILLCELL_220_512 ();
 FILLCELL_X32 FILLCELL_220_544 ();
 FILLCELL_X32 FILLCELL_220_576 ();
 FILLCELL_X32 FILLCELL_220_608 ();
 FILLCELL_X32 FILLCELL_220_640 ();
 FILLCELL_X32 FILLCELL_220_672 ();
 FILLCELL_X32 FILLCELL_220_704 ();
 FILLCELL_X32 FILLCELL_220_736 ();
 FILLCELL_X32 FILLCELL_220_768 ();
 FILLCELL_X32 FILLCELL_220_800 ();
 FILLCELL_X32 FILLCELL_220_832 ();
 FILLCELL_X32 FILLCELL_220_864 ();
 FILLCELL_X32 FILLCELL_220_896 ();
 FILLCELL_X32 FILLCELL_220_928 ();
 FILLCELL_X32 FILLCELL_220_960 ();
 FILLCELL_X32 FILLCELL_220_992 ();
 FILLCELL_X32 FILLCELL_220_1024 ();
 FILLCELL_X32 FILLCELL_220_1056 ();
 FILLCELL_X32 FILLCELL_220_1088 ();
 FILLCELL_X32 FILLCELL_220_1120 ();
 FILLCELL_X32 FILLCELL_220_1152 ();
 FILLCELL_X32 FILLCELL_220_1184 ();
 FILLCELL_X32 FILLCELL_220_1216 ();
 FILLCELL_X32 FILLCELL_220_1248 ();
 FILLCELL_X32 FILLCELL_220_1280 ();
 FILLCELL_X32 FILLCELL_220_1312 ();
 FILLCELL_X32 FILLCELL_220_1344 ();
 FILLCELL_X32 FILLCELL_220_1376 ();
 FILLCELL_X32 FILLCELL_220_1408 ();
 FILLCELL_X32 FILLCELL_220_1440 ();
 FILLCELL_X32 FILLCELL_220_1472 ();
 FILLCELL_X32 FILLCELL_220_1504 ();
 FILLCELL_X32 FILLCELL_220_1536 ();
 FILLCELL_X32 FILLCELL_220_1568 ();
 FILLCELL_X32 FILLCELL_220_1600 ();
 FILLCELL_X32 FILLCELL_220_1632 ();
 FILLCELL_X32 FILLCELL_220_1664 ();
 FILLCELL_X32 FILLCELL_220_1696 ();
 FILLCELL_X32 FILLCELL_220_1728 ();
 FILLCELL_X32 FILLCELL_220_1760 ();
 FILLCELL_X32 FILLCELL_220_1792 ();
 FILLCELL_X32 FILLCELL_220_1824 ();
 FILLCELL_X32 FILLCELL_220_1856 ();
 FILLCELL_X8 FILLCELL_220_1888 ();
 FILLCELL_X1 FILLCELL_220_1896 ();
 FILLCELL_X32 FILLCELL_221_0 ();
 FILLCELL_X32 FILLCELL_221_32 ();
 FILLCELL_X32 FILLCELL_221_64 ();
 FILLCELL_X32 FILLCELL_221_96 ();
 FILLCELL_X32 FILLCELL_221_128 ();
 FILLCELL_X32 FILLCELL_221_160 ();
 FILLCELL_X32 FILLCELL_221_192 ();
 FILLCELL_X32 FILLCELL_221_224 ();
 FILLCELL_X32 FILLCELL_221_256 ();
 FILLCELL_X32 FILLCELL_221_288 ();
 FILLCELL_X32 FILLCELL_221_320 ();
 FILLCELL_X32 FILLCELL_221_352 ();
 FILLCELL_X32 FILLCELL_221_384 ();
 FILLCELL_X32 FILLCELL_221_416 ();
 FILLCELL_X32 FILLCELL_221_448 ();
 FILLCELL_X32 FILLCELL_221_480 ();
 FILLCELL_X32 FILLCELL_221_512 ();
 FILLCELL_X32 FILLCELL_221_544 ();
 FILLCELL_X32 FILLCELL_221_576 ();
 FILLCELL_X32 FILLCELL_221_608 ();
 FILLCELL_X32 FILLCELL_221_640 ();
 FILLCELL_X32 FILLCELL_221_672 ();
 FILLCELL_X32 FILLCELL_221_704 ();
 FILLCELL_X32 FILLCELL_221_736 ();
 FILLCELL_X32 FILLCELL_221_768 ();
 FILLCELL_X32 FILLCELL_221_800 ();
 FILLCELL_X32 FILLCELL_221_832 ();
 FILLCELL_X32 FILLCELL_221_864 ();
 FILLCELL_X32 FILLCELL_221_896 ();
 FILLCELL_X32 FILLCELL_221_928 ();
 FILLCELL_X32 FILLCELL_221_960 ();
 FILLCELL_X32 FILLCELL_221_992 ();
 FILLCELL_X32 FILLCELL_221_1024 ();
 FILLCELL_X32 FILLCELL_221_1056 ();
 FILLCELL_X32 FILLCELL_221_1088 ();
 FILLCELL_X32 FILLCELL_221_1120 ();
 FILLCELL_X32 FILLCELL_221_1152 ();
 FILLCELL_X32 FILLCELL_221_1184 ();
 FILLCELL_X32 FILLCELL_221_1216 ();
 FILLCELL_X32 FILLCELL_221_1248 ();
 FILLCELL_X32 FILLCELL_221_1280 ();
 FILLCELL_X32 FILLCELL_221_1312 ();
 FILLCELL_X32 FILLCELL_221_1344 ();
 FILLCELL_X32 FILLCELL_221_1376 ();
 FILLCELL_X32 FILLCELL_221_1408 ();
 FILLCELL_X32 FILLCELL_221_1440 ();
 FILLCELL_X32 FILLCELL_221_1472 ();
 FILLCELL_X32 FILLCELL_221_1504 ();
 FILLCELL_X32 FILLCELL_221_1536 ();
 FILLCELL_X32 FILLCELL_221_1568 ();
 FILLCELL_X32 FILLCELL_221_1600 ();
 FILLCELL_X32 FILLCELL_221_1632 ();
 FILLCELL_X32 FILLCELL_221_1664 ();
 FILLCELL_X32 FILLCELL_221_1696 ();
 FILLCELL_X32 FILLCELL_221_1728 ();
 FILLCELL_X32 FILLCELL_221_1760 ();
 FILLCELL_X32 FILLCELL_221_1792 ();
 FILLCELL_X32 FILLCELL_221_1824 ();
 FILLCELL_X32 FILLCELL_221_1856 ();
 FILLCELL_X8 FILLCELL_221_1888 ();
 FILLCELL_X1 FILLCELL_221_1896 ();
 FILLCELL_X32 FILLCELL_222_0 ();
 FILLCELL_X32 FILLCELL_222_32 ();
 FILLCELL_X32 FILLCELL_222_64 ();
 FILLCELL_X32 FILLCELL_222_96 ();
 FILLCELL_X32 FILLCELL_222_128 ();
 FILLCELL_X32 FILLCELL_222_160 ();
 FILLCELL_X32 FILLCELL_222_192 ();
 FILLCELL_X32 FILLCELL_222_224 ();
 FILLCELL_X32 FILLCELL_222_256 ();
 FILLCELL_X32 FILLCELL_222_288 ();
 FILLCELL_X32 FILLCELL_222_320 ();
 FILLCELL_X32 FILLCELL_222_352 ();
 FILLCELL_X32 FILLCELL_222_384 ();
 FILLCELL_X32 FILLCELL_222_416 ();
 FILLCELL_X32 FILLCELL_222_448 ();
 FILLCELL_X32 FILLCELL_222_480 ();
 FILLCELL_X32 FILLCELL_222_512 ();
 FILLCELL_X32 FILLCELL_222_544 ();
 FILLCELL_X32 FILLCELL_222_576 ();
 FILLCELL_X32 FILLCELL_222_608 ();
 FILLCELL_X32 FILLCELL_222_640 ();
 FILLCELL_X32 FILLCELL_222_672 ();
 FILLCELL_X32 FILLCELL_222_704 ();
 FILLCELL_X32 FILLCELL_222_736 ();
 FILLCELL_X32 FILLCELL_222_768 ();
 FILLCELL_X32 FILLCELL_222_800 ();
 FILLCELL_X32 FILLCELL_222_832 ();
 FILLCELL_X32 FILLCELL_222_864 ();
 FILLCELL_X32 FILLCELL_222_896 ();
 FILLCELL_X32 FILLCELL_222_928 ();
 FILLCELL_X32 FILLCELL_222_960 ();
 FILLCELL_X32 FILLCELL_222_992 ();
 FILLCELL_X32 FILLCELL_222_1024 ();
 FILLCELL_X32 FILLCELL_222_1056 ();
 FILLCELL_X32 FILLCELL_222_1088 ();
 FILLCELL_X32 FILLCELL_222_1120 ();
 FILLCELL_X32 FILLCELL_222_1152 ();
 FILLCELL_X32 FILLCELL_222_1184 ();
 FILLCELL_X32 FILLCELL_222_1216 ();
 FILLCELL_X32 FILLCELL_222_1248 ();
 FILLCELL_X32 FILLCELL_222_1280 ();
 FILLCELL_X32 FILLCELL_222_1312 ();
 FILLCELL_X32 FILLCELL_222_1344 ();
 FILLCELL_X32 FILLCELL_222_1376 ();
 FILLCELL_X32 FILLCELL_222_1408 ();
 FILLCELL_X32 FILLCELL_222_1440 ();
 FILLCELL_X32 FILLCELL_222_1472 ();
 FILLCELL_X32 FILLCELL_222_1504 ();
 FILLCELL_X32 FILLCELL_222_1536 ();
 FILLCELL_X32 FILLCELL_222_1568 ();
 FILLCELL_X32 FILLCELL_222_1600 ();
 FILLCELL_X32 FILLCELL_222_1632 ();
 FILLCELL_X32 FILLCELL_222_1664 ();
 FILLCELL_X32 FILLCELL_222_1696 ();
 FILLCELL_X32 FILLCELL_222_1728 ();
 FILLCELL_X32 FILLCELL_222_1760 ();
 FILLCELL_X32 FILLCELL_222_1792 ();
 FILLCELL_X32 FILLCELL_222_1824 ();
 FILLCELL_X32 FILLCELL_222_1856 ();
 FILLCELL_X8 FILLCELL_222_1888 ();
 FILLCELL_X1 FILLCELL_222_1896 ();
 FILLCELL_X32 FILLCELL_223_0 ();
 FILLCELL_X32 FILLCELL_223_32 ();
 FILLCELL_X32 FILLCELL_223_64 ();
 FILLCELL_X32 FILLCELL_223_96 ();
 FILLCELL_X32 FILLCELL_223_128 ();
 FILLCELL_X32 FILLCELL_223_160 ();
 FILLCELL_X32 FILLCELL_223_192 ();
 FILLCELL_X32 FILLCELL_223_224 ();
 FILLCELL_X32 FILLCELL_223_256 ();
 FILLCELL_X32 FILLCELL_223_288 ();
 FILLCELL_X32 FILLCELL_223_320 ();
 FILLCELL_X32 FILLCELL_223_352 ();
 FILLCELL_X32 FILLCELL_223_384 ();
 FILLCELL_X32 FILLCELL_223_416 ();
 FILLCELL_X32 FILLCELL_223_448 ();
 FILLCELL_X32 FILLCELL_223_480 ();
 FILLCELL_X32 FILLCELL_223_512 ();
 FILLCELL_X32 FILLCELL_223_544 ();
 FILLCELL_X32 FILLCELL_223_576 ();
 FILLCELL_X32 FILLCELL_223_608 ();
 FILLCELL_X32 FILLCELL_223_640 ();
 FILLCELL_X32 FILLCELL_223_672 ();
 FILLCELL_X32 FILLCELL_223_704 ();
 FILLCELL_X32 FILLCELL_223_736 ();
 FILLCELL_X32 FILLCELL_223_768 ();
 FILLCELL_X32 FILLCELL_223_800 ();
 FILLCELL_X32 FILLCELL_223_832 ();
 FILLCELL_X32 FILLCELL_223_864 ();
 FILLCELL_X32 FILLCELL_223_896 ();
 FILLCELL_X32 FILLCELL_223_928 ();
 FILLCELL_X32 FILLCELL_223_960 ();
 FILLCELL_X32 FILLCELL_223_992 ();
 FILLCELL_X32 FILLCELL_223_1024 ();
 FILLCELL_X32 FILLCELL_223_1056 ();
 FILLCELL_X32 FILLCELL_223_1088 ();
 FILLCELL_X32 FILLCELL_223_1120 ();
 FILLCELL_X32 FILLCELL_223_1152 ();
 FILLCELL_X32 FILLCELL_223_1184 ();
 FILLCELL_X32 FILLCELL_223_1216 ();
 FILLCELL_X32 FILLCELL_223_1248 ();
 FILLCELL_X32 FILLCELL_223_1280 ();
 FILLCELL_X32 FILLCELL_223_1312 ();
 FILLCELL_X32 FILLCELL_223_1344 ();
 FILLCELL_X32 FILLCELL_223_1376 ();
 FILLCELL_X32 FILLCELL_223_1408 ();
 FILLCELL_X32 FILLCELL_223_1440 ();
 FILLCELL_X32 FILLCELL_223_1472 ();
 FILLCELL_X32 FILLCELL_223_1504 ();
 FILLCELL_X32 FILLCELL_223_1536 ();
 FILLCELL_X32 FILLCELL_223_1568 ();
 FILLCELL_X32 FILLCELL_223_1600 ();
 FILLCELL_X32 FILLCELL_223_1632 ();
 FILLCELL_X32 FILLCELL_223_1664 ();
 FILLCELL_X32 FILLCELL_223_1696 ();
 FILLCELL_X32 FILLCELL_223_1728 ();
 FILLCELL_X32 FILLCELL_223_1760 ();
 FILLCELL_X32 FILLCELL_223_1792 ();
 FILLCELL_X32 FILLCELL_223_1824 ();
 FILLCELL_X32 FILLCELL_223_1856 ();
 FILLCELL_X8 FILLCELL_223_1888 ();
 FILLCELL_X1 FILLCELL_223_1896 ();
 FILLCELL_X32 FILLCELL_224_0 ();
 FILLCELL_X32 FILLCELL_224_32 ();
 FILLCELL_X32 FILLCELL_224_64 ();
 FILLCELL_X32 FILLCELL_224_96 ();
 FILLCELL_X32 FILLCELL_224_128 ();
 FILLCELL_X32 FILLCELL_224_160 ();
 FILLCELL_X32 FILLCELL_224_192 ();
 FILLCELL_X32 FILLCELL_224_224 ();
 FILLCELL_X32 FILLCELL_224_256 ();
 FILLCELL_X32 FILLCELL_224_288 ();
 FILLCELL_X32 FILLCELL_224_320 ();
 FILLCELL_X32 FILLCELL_224_352 ();
 FILLCELL_X32 FILLCELL_224_384 ();
 FILLCELL_X32 FILLCELL_224_416 ();
 FILLCELL_X32 FILLCELL_224_448 ();
 FILLCELL_X32 FILLCELL_224_480 ();
 FILLCELL_X32 FILLCELL_224_512 ();
 FILLCELL_X32 FILLCELL_224_544 ();
 FILLCELL_X32 FILLCELL_224_576 ();
 FILLCELL_X32 FILLCELL_224_608 ();
 FILLCELL_X32 FILLCELL_224_640 ();
 FILLCELL_X32 FILLCELL_224_672 ();
 FILLCELL_X32 FILLCELL_224_704 ();
 FILLCELL_X32 FILLCELL_224_736 ();
 FILLCELL_X32 FILLCELL_224_768 ();
 FILLCELL_X32 FILLCELL_224_800 ();
 FILLCELL_X32 FILLCELL_224_832 ();
 FILLCELL_X32 FILLCELL_224_864 ();
 FILLCELL_X32 FILLCELL_224_896 ();
 FILLCELL_X32 FILLCELL_224_928 ();
 FILLCELL_X32 FILLCELL_224_960 ();
 FILLCELL_X32 FILLCELL_224_992 ();
 FILLCELL_X32 FILLCELL_224_1024 ();
 FILLCELL_X32 FILLCELL_224_1056 ();
 FILLCELL_X32 FILLCELL_224_1088 ();
 FILLCELL_X32 FILLCELL_224_1120 ();
 FILLCELL_X32 FILLCELL_224_1152 ();
 FILLCELL_X32 FILLCELL_224_1184 ();
 FILLCELL_X32 FILLCELL_224_1216 ();
 FILLCELL_X32 FILLCELL_224_1248 ();
 FILLCELL_X32 FILLCELL_224_1280 ();
 FILLCELL_X32 FILLCELL_224_1312 ();
 FILLCELL_X32 FILLCELL_224_1344 ();
 FILLCELL_X32 FILLCELL_224_1376 ();
 FILLCELL_X32 FILLCELL_224_1408 ();
 FILLCELL_X32 FILLCELL_224_1440 ();
 FILLCELL_X32 FILLCELL_224_1472 ();
 FILLCELL_X32 FILLCELL_224_1504 ();
 FILLCELL_X32 FILLCELL_224_1536 ();
 FILLCELL_X32 FILLCELL_224_1568 ();
 FILLCELL_X32 FILLCELL_224_1600 ();
 FILLCELL_X32 FILLCELL_224_1632 ();
 FILLCELL_X32 FILLCELL_224_1664 ();
 FILLCELL_X32 FILLCELL_224_1696 ();
 FILLCELL_X32 FILLCELL_224_1728 ();
 FILLCELL_X32 FILLCELL_224_1760 ();
 FILLCELL_X32 FILLCELL_224_1792 ();
 FILLCELL_X32 FILLCELL_224_1824 ();
 FILLCELL_X32 FILLCELL_224_1856 ();
 FILLCELL_X8 FILLCELL_224_1888 ();
 FILLCELL_X1 FILLCELL_224_1896 ();
 FILLCELL_X32 FILLCELL_225_0 ();
 FILLCELL_X32 FILLCELL_225_32 ();
 FILLCELL_X32 FILLCELL_225_64 ();
 FILLCELL_X32 FILLCELL_225_96 ();
 FILLCELL_X32 FILLCELL_225_128 ();
 FILLCELL_X32 FILLCELL_225_160 ();
 FILLCELL_X32 FILLCELL_225_192 ();
 FILLCELL_X32 FILLCELL_225_224 ();
 FILLCELL_X32 FILLCELL_225_256 ();
 FILLCELL_X32 FILLCELL_225_288 ();
 FILLCELL_X32 FILLCELL_225_320 ();
 FILLCELL_X32 FILLCELL_225_352 ();
 FILLCELL_X32 FILLCELL_225_384 ();
 FILLCELL_X32 FILLCELL_225_416 ();
 FILLCELL_X32 FILLCELL_225_448 ();
 FILLCELL_X32 FILLCELL_225_480 ();
 FILLCELL_X32 FILLCELL_225_512 ();
 FILLCELL_X32 FILLCELL_225_544 ();
 FILLCELL_X32 FILLCELL_225_576 ();
 FILLCELL_X32 FILLCELL_225_608 ();
 FILLCELL_X32 FILLCELL_225_640 ();
 FILLCELL_X32 FILLCELL_225_672 ();
 FILLCELL_X32 FILLCELL_225_704 ();
 FILLCELL_X32 FILLCELL_225_736 ();
 FILLCELL_X32 FILLCELL_225_768 ();
 FILLCELL_X32 FILLCELL_225_800 ();
 FILLCELL_X32 FILLCELL_225_832 ();
 FILLCELL_X32 FILLCELL_225_864 ();
 FILLCELL_X32 FILLCELL_225_896 ();
 FILLCELL_X32 FILLCELL_225_928 ();
 FILLCELL_X32 FILLCELL_225_960 ();
 FILLCELL_X32 FILLCELL_225_992 ();
 FILLCELL_X32 FILLCELL_225_1024 ();
 FILLCELL_X32 FILLCELL_225_1056 ();
 FILLCELL_X32 FILLCELL_225_1088 ();
 FILLCELL_X32 FILLCELL_225_1120 ();
 FILLCELL_X32 FILLCELL_225_1152 ();
 FILLCELL_X32 FILLCELL_225_1184 ();
 FILLCELL_X32 FILLCELL_225_1216 ();
 FILLCELL_X32 FILLCELL_225_1248 ();
 FILLCELL_X32 FILLCELL_225_1280 ();
 FILLCELL_X32 FILLCELL_225_1312 ();
 FILLCELL_X32 FILLCELL_225_1344 ();
 FILLCELL_X32 FILLCELL_225_1376 ();
 FILLCELL_X32 FILLCELL_225_1408 ();
 FILLCELL_X32 FILLCELL_225_1440 ();
 FILLCELL_X32 FILLCELL_225_1472 ();
 FILLCELL_X32 FILLCELL_225_1504 ();
 FILLCELL_X32 FILLCELL_225_1536 ();
 FILLCELL_X32 FILLCELL_225_1568 ();
 FILLCELL_X32 FILLCELL_225_1600 ();
 FILLCELL_X32 FILLCELL_225_1632 ();
 FILLCELL_X32 FILLCELL_225_1664 ();
 FILLCELL_X32 FILLCELL_225_1696 ();
 FILLCELL_X32 FILLCELL_225_1728 ();
 FILLCELL_X32 FILLCELL_225_1760 ();
 FILLCELL_X32 FILLCELL_225_1792 ();
 FILLCELL_X32 FILLCELL_225_1824 ();
 FILLCELL_X32 FILLCELL_225_1856 ();
 FILLCELL_X8 FILLCELL_225_1888 ();
 FILLCELL_X1 FILLCELL_225_1896 ();
 FILLCELL_X32 FILLCELL_226_0 ();
 FILLCELL_X32 FILLCELL_226_32 ();
 FILLCELL_X32 FILLCELL_226_64 ();
 FILLCELL_X32 FILLCELL_226_96 ();
 FILLCELL_X32 FILLCELL_226_128 ();
 FILLCELL_X32 FILLCELL_226_160 ();
 FILLCELL_X32 FILLCELL_226_192 ();
 FILLCELL_X32 FILLCELL_226_224 ();
 FILLCELL_X32 FILLCELL_226_256 ();
 FILLCELL_X32 FILLCELL_226_288 ();
 FILLCELL_X32 FILLCELL_226_320 ();
 FILLCELL_X32 FILLCELL_226_352 ();
 FILLCELL_X32 FILLCELL_226_384 ();
 FILLCELL_X32 FILLCELL_226_416 ();
 FILLCELL_X32 FILLCELL_226_448 ();
 FILLCELL_X32 FILLCELL_226_480 ();
 FILLCELL_X32 FILLCELL_226_512 ();
 FILLCELL_X32 FILLCELL_226_544 ();
 FILLCELL_X32 FILLCELL_226_576 ();
 FILLCELL_X32 FILLCELL_226_608 ();
 FILLCELL_X32 FILLCELL_226_640 ();
 FILLCELL_X32 FILLCELL_226_672 ();
 FILLCELL_X32 FILLCELL_226_704 ();
 FILLCELL_X32 FILLCELL_226_736 ();
 FILLCELL_X32 FILLCELL_226_768 ();
 FILLCELL_X32 FILLCELL_226_800 ();
 FILLCELL_X32 FILLCELL_226_832 ();
 FILLCELL_X32 FILLCELL_226_864 ();
 FILLCELL_X32 FILLCELL_226_896 ();
 FILLCELL_X32 FILLCELL_226_928 ();
 FILLCELL_X32 FILLCELL_226_960 ();
 FILLCELL_X32 FILLCELL_226_992 ();
 FILLCELL_X32 FILLCELL_226_1024 ();
 FILLCELL_X32 FILLCELL_226_1056 ();
 FILLCELL_X32 FILLCELL_226_1088 ();
 FILLCELL_X32 FILLCELL_226_1120 ();
 FILLCELL_X32 FILLCELL_226_1152 ();
 FILLCELL_X32 FILLCELL_226_1184 ();
 FILLCELL_X32 FILLCELL_226_1216 ();
 FILLCELL_X32 FILLCELL_226_1248 ();
 FILLCELL_X32 FILLCELL_226_1280 ();
 FILLCELL_X32 FILLCELL_226_1312 ();
 FILLCELL_X32 FILLCELL_226_1344 ();
 FILLCELL_X32 FILLCELL_226_1376 ();
 FILLCELL_X32 FILLCELL_226_1408 ();
 FILLCELL_X32 FILLCELL_226_1440 ();
 FILLCELL_X32 FILLCELL_226_1472 ();
 FILLCELL_X32 FILLCELL_226_1504 ();
 FILLCELL_X32 FILLCELL_226_1536 ();
 FILLCELL_X32 FILLCELL_226_1568 ();
 FILLCELL_X32 FILLCELL_226_1600 ();
 FILLCELL_X32 FILLCELL_226_1632 ();
 FILLCELL_X32 FILLCELL_226_1664 ();
 FILLCELL_X32 FILLCELL_226_1696 ();
 FILLCELL_X32 FILLCELL_226_1728 ();
 FILLCELL_X32 FILLCELL_226_1760 ();
 FILLCELL_X32 FILLCELL_226_1792 ();
 FILLCELL_X32 FILLCELL_226_1824 ();
 FILLCELL_X32 FILLCELL_226_1856 ();
 FILLCELL_X8 FILLCELL_226_1888 ();
 FILLCELL_X1 FILLCELL_226_1896 ();
 FILLCELL_X32 FILLCELL_227_0 ();
 FILLCELL_X32 FILLCELL_227_32 ();
 FILLCELL_X32 FILLCELL_227_64 ();
 FILLCELL_X32 FILLCELL_227_96 ();
 FILLCELL_X32 FILLCELL_227_128 ();
 FILLCELL_X32 FILLCELL_227_160 ();
 FILLCELL_X32 FILLCELL_227_192 ();
 FILLCELL_X32 FILLCELL_227_224 ();
 FILLCELL_X32 FILLCELL_227_256 ();
 FILLCELL_X32 FILLCELL_227_288 ();
 FILLCELL_X32 FILLCELL_227_320 ();
 FILLCELL_X32 FILLCELL_227_352 ();
 FILLCELL_X32 FILLCELL_227_384 ();
 FILLCELL_X32 FILLCELL_227_416 ();
 FILLCELL_X32 FILLCELL_227_448 ();
 FILLCELL_X32 FILLCELL_227_480 ();
 FILLCELL_X32 FILLCELL_227_512 ();
 FILLCELL_X32 FILLCELL_227_544 ();
 FILLCELL_X32 FILLCELL_227_576 ();
 FILLCELL_X32 FILLCELL_227_608 ();
 FILLCELL_X32 FILLCELL_227_640 ();
 FILLCELL_X32 FILLCELL_227_672 ();
 FILLCELL_X32 FILLCELL_227_704 ();
 FILLCELL_X32 FILLCELL_227_736 ();
 FILLCELL_X32 FILLCELL_227_768 ();
 FILLCELL_X32 FILLCELL_227_800 ();
 FILLCELL_X32 FILLCELL_227_832 ();
 FILLCELL_X32 FILLCELL_227_864 ();
 FILLCELL_X32 FILLCELL_227_896 ();
 FILLCELL_X32 FILLCELL_227_928 ();
 FILLCELL_X32 FILLCELL_227_960 ();
 FILLCELL_X32 FILLCELL_227_992 ();
 FILLCELL_X32 FILLCELL_227_1024 ();
 FILLCELL_X32 FILLCELL_227_1056 ();
 FILLCELL_X32 FILLCELL_227_1088 ();
 FILLCELL_X32 FILLCELL_227_1120 ();
 FILLCELL_X32 FILLCELL_227_1152 ();
 FILLCELL_X32 FILLCELL_227_1184 ();
 FILLCELL_X32 FILLCELL_227_1216 ();
 FILLCELL_X32 FILLCELL_227_1248 ();
 FILLCELL_X32 FILLCELL_227_1280 ();
 FILLCELL_X32 FILLCELL_227_1312 ();
 FILLCELL_X32 FILLCELL_227_1344 ();
 FILLCELL_X32 FILLCELL_227_1376 ();
 FILLCELL_X32 FILLCELL_227_1408 ();
 FILLCELL_X32 FILLCELL_227_1440 ();
 FILLCELL_X32 FILLCELL_227_1472 ();
 FILLCELL_X32 FILLCELL_227_1504 ();
 FILLCELL_X32 FILLCELL_227_1536 ();
 FILLCELL_X32 FILLCELL_227_1568 ();
 FILLCELL_X32 FILLCELL_227_1600 ();
 FILLCELL_X32 FILLCELL_227_1632 ();
 FILLCELL_X32 FILLCELL_227_1664 ();
 FILLCELL_X32 FILLCELL_227_1696 ();
 FILLCELL_X32 FILLCELL_227_1728 ();
 FILLCELL_X32 FILLCELL_227_1760 ();
 FILLCELL_X32 FILLCELL_227_1792 ();
 FILLCELL_X32 FILLCELL_227_1824 ();
 FILLCELL_X32 FILLCELL_227_1856 ();
 FILLCELL_X8 FILLCELL_227_1888 ();
 FILLCELL_X1 FILLCELL_227_1896 ();
 FILLCELL_X32 FILLCELL_228_0 ();
 FILLCELL_X32 FILLCELL_228_32 ();
 FILLCELL_X32 FILLCELL_228_64 ();
 FILLCELL_X32 FILLCELL_228_96 ();
 FILLCELL_X32 FILLCELL_228_128 ();
 FILLCELL_X32 FILLCELL_228_160 ();
 FILLCELL_X32 FILLCELL_228_192 ();
 FILLCELL_X32 FILLCELL_228_224 ();
 FILLCELL_X32 FILLCELL_228_256 ();
 FILLCELL_X32 FILLCELL_228_288 ();
 FILLCELL_X32 FILLCELL_228_320 ();
 FILLCELL_X32 FILLCELL_228_352 ();
 FILLCELL_X32 FILLCELL_228_384 ();
 FILLCELL_X32 FILLCELL_228_416 ();
 FILLCELL_X32 FILLCELL_228_448 ();
 FILLCELL_X32 FILLCELL_228_480 ();
 FILLCELL_X32 FILLCELL_228_512 ();
 FILLCELL_X32 FILLCELL_228_544 ();
 FILLCELL_X32 FILLCELL_228_576 ();
 FILLCELL_X32 FILLCELL_228_608 ();
 FILLCELL_X32 FILLCELL_228_640 ();
 FILLCELL_X32 FILLCELL_228_672 ();
 FILLCELL_X32 FILLCELL_228_704 ();
 FILLCELL_X32 FILLCELL_228_736 ();
 FILLCELL_X32 FILLCELL_228_768 ();
 FILLCELL_X32 FILLCELL_228_800 ();
 FILLCELL_X32 FILLCELL_228_832 ();
 FILLCELL_X32 FILLCELL_228_864 ();
 FILLCELL_X32 FILLCELL_228_896 ();
 FILLCELL_X32 FILLCELL_228_928 ();
 FILLCELL_X32 FILLCELL_228_960 ();
 FILLCELL_X32 FILLCELL_228_992 ();
 FILLCELL_X32 FILLCELL_228_1024 ();
 FILLCELL_X32 FILLCELL_228_1056 ();
 FILLCELL_X32 FILLCELL_228_1088 ();
 FILLCELL_X32 FILLCELL_228_1120 ();
 FILLCELL_X32 FILLCELL_228_1152 ();
 FILLCELL_X32 FILLCELL_228_1184 ();
 FILLCELL_X32 FILLCELL_228_1216 ();
 FILLCELL_X32 FILLCELL_228_1248 ();
 FILLCELL_X32 FILLCELL_228_1280 ();
 FILLCELL_X32 FILLCELL_228_1312 ();
 FILLCELL_X32 FILLCELL_228_1344 ();
 FILLCELL_X32 FILLCELL_228_1376 ();
 FILLCELL_X32 FILLCELL_228_1408 ();
 FILLCELL_X32 FILLCELL_228_1440 ();
 FILLCELL_X32 FILLCELL_228_1472 ();
 FILLCELL_X32 FILLCELL_228_1504 ();
 FILLCELL_X32 FILLCELL_228_1536 ();
 FILLCELL_X32 FILLCELL_228_1568 ();
 FILLCELL_X32 FILLCELL_228_1600 ();
 FILLCELL_X32 FILLCELL_228_1632 ();
 FILLCELL_X32 FILLCELL_228_1664 ();
 FILLCELL_X32 FILLCELL_228_1696 ();
 FILLCELL_X32 FILLCELL_228_1728 ();
 FILLCELL_X32 FILLCELL_228_1760 ();
 FILLCELL_X32 FILLCELL_228_1792 ();
 FILLCELL_X32 FILLCELL_228_1824 ();
 FILLCELL_X32 FILLCELL_228_1856 ();
 FILLCELL_X8 FILLCELL_228_1888 ();
 FILLCELL_X1 FILLCELL_228_1896 ();
 FILLCELL_X32 FILLCELL_229_0 ();
 FILLCELL_X32 FILLCELL_229_32 ();
 FILLCELL_X32 FILLCELL_229_64 ();
 FILLCELL_X32 FILLCELL_229_96 ();
 FILLCELL_X32 FILLCELL_229_128 ();
 FILLCELL_X32 FILLCELL_229_160 ();
 FILLCELL_X32 FILLCELL_229_192 ();
 FILLCELL_X32 FILLCELL_229_224 ();
 FILLCELL_X32 FILLCELL_229_256 ();
 FILLCELL_X32 FILLCELL_229_288 ();
 FILLCELL_X32 FILLCELL_229_320 ();
 FILLCELL_X32 FILLCELL_229_352 ();
 FILLCELL_X32 FILLCELL_229_384 ();
 FILLCELL_X32 FILLCELL_229_416 ();
 FILLCELL_X32 FILLCELL_229_448 ();
 FILLCELL_X32 FILLCELL_229_480 ();
 FILLCELL_X32 FILLCELL_229_512 ();
 FILLCELL_X32 FILLCELL_229_544 ();
 FILLCELL_X32 FILLCELL_229_576 ();
 FILLCELL_X32 FILLCELL_229_608 ();
 FILLCELL_X32 FILLCELL_229_640 ();
 FILLCELL_X32 FILLCELL_229_672 ();
 FILLCELL_X32 FILLCELL_229_704 ();
 FILLCELL_X32 FILLCELL_229_736 ();
 FILLCELL_X32 FILLCELL_229_768 ();
 FILLCELL_X32 FILLCELL_229_800 ();
 FILLCELL_X32 FILLCELL_229_832 ();
 FILLCELL_X32 FILLCELL_229_864 ();
 FILLCELL_X32 FILLCELL_229_896 ();
 FILLCELL_X32 FILLCELL_229_928 ();
 FILLCELL_X32 FILLCELL_229_960 ();
 FILLCELL_X32 FILLCELL_229_992 ();
 FILLCELL_X32 FILLCELL_229_1024 ();
 FILLCELL_X32 FILLCELL_229_1056 ();
 FILLCELL_X32 FILLCELL_229_1088 ();
 FILLCELL_X32 FILLCELL_229_1120 ();
 FILLCELL_X32 FILLCELL_229_1152 ();
 FILLCELL_X32 FILLCELL_229_1184 ();
 FILLCELL_X32 FILLCELL_229_1216 ();
 FILLCELL_X32 FILLCELL_229_1248 ();
 FILLCELL_X32 FILLCELL_229_1280 ();
 FILLCELL_X32 FILLCELL_229_1312 ();
 FILLCELL_X32 FILLCELL_229_1344 ();
 FILLCELL_X32 FILLCELL_229_1376 ();
 FILLCELL_X32 FILLCELL_229_1408 ();
 FILLCELL_X32 FILLCELL_229_1440 ();
 FILLCELL_X32 FILLCELL_229_1472 ();
 FILLCELL_X32 FILLCELL_229_1504 ();
 FILLCELL_X32 FILLCELL_229_1536 ();
 FILLCELL_X32 FILLCELL_229_1568 ();
 FILLCELL_X32 FILLCELL_229_1600 ();
 FILLCELL_X32 FILLCELL_229_1632 ();
 FILLCELL_X32 FILLCELL_229_1664 ();
 FILLCELL_X32 FILLCELL_229_1696 ();
 FILLCELL_X32 FILLCELL_229_1728 ();
 FILLCELL_X32 FILLCELL_229_1760 ();
 FILLCELL_X32 FILLCELL_229_1792 ();
 FILLCELL_X32 FILLCELL_229_1824 ();
 FILLCELL_X32 FILLCELL_229_1856 ();
 FILLCELL_X8 FILLCELL_229_1888 ();
 FILLCELL_X1 FILLCELL_229_1896 ();
 FILLCELL_X32 FILLCELL_230_0 ();
 FILLCELL_X32 FILLCELL_230_32 ();
 FILLCELL_X32 FILLCELL_230_64 ();
 FILLCELL_X32 FILLCELL_230_96 ();
 FILLCELL_X32 FILLCELL_230_128 ();
 FILLCELL_X32 FILLCELL_230_160 ();
 FILLCELL_X32 FILLCELL_230_192 ();
 FILLCELL_X32 FILLCELL_230_224 ();
 FILLCELL_X32 FILLCELL_230_256 ();
 FILLCELL_X32 FILLCELL_230_288 ();
 FILLCELL_X32 FILLCELL_230_320 ();
 FILLCELL_X32 FILLCELL_230_352 ();
 FILLCELL_X32 FILLCELL_230_384 ();
 FILLCELL_X32 FILLCELL_230_416 ();
 FILLCELL_X32 FILLCELL_230_448 ();
 FILLCELL_X32 FILLCELL_230_480 ();
 FILLCELL_X32 FILLCELL_230_512 ();
 FILLCELL_X32 FILLCELL_230_544 ();
 FILLCELL_X32 FILLCELL_230_576 ();
 FILLCELL_X32 FILLCELL_230_608 ();
 FILLCELL_X32 FILLCELL_230_640 ();
 FILLCELL_X32 FILLCELL_230_672 ();
 FILLCELL_X32 FILLCELL_230_704 ();
 FILLCELL_X32 FILLCELL_230_736 ();
 FILLCELL_X32 FILLCELL_230_768 ();
 FILLCELL_X32 FILLCELL_230_800 ();
 FILLCELL_X32 FILLCELL_230_832 ();
 FILLCELL_X32 FILLCELL_230_864 ();
 FILLCELL_X32 FILLCELL_230_896 ();
 FILLCELL_X32 FILLCELL_230_928 ();
 FILLCELL_X32 FILLCELL_230_960 ();
 FILLCELL_X32 FILLCELL_230_992 ();
 FILLCELL_X32 FILLCELL_230_1024 ();
 FILLCELL_X32 FILLCELL_230_1056 ();
 FILLCELL_X32 FILLCELL_230_1088 ();
 FILLCELL_X32 FILLCELL_230_1120 ();
 FILLCELL_X32 FILLCELL_230_1152 ();
 FILLCELL_X32 FILLCELL_230_1184 ();
 FILLCELL_X32 FILLCELL_230_1216 ();
 FILLCELL_X32 FILLCELL_230_1248 ();
 FILLCELL_X32 FILLCELL_230_1280 ();
 FILLCELL_X32 FILLCELL_230_1312 ();
 FILLCELL_X32 FILLCELL_230_1344 ();
 FILLCELL_X32 FILLCELL_230_1376 ();
 FILLCELL_X32 FILLCELL_230_1408 ();
 FILLCELL_X32 FILLCELL_230_1440 ();
 FILLCELL_X32 FILLCELL_230_1472 ();
 FILLCELL_X32 FILLCELL_230_1504 ();
 FILLCELL_X32 FILLCELL_230_1536 ();
 FILLCELL_X32 FILLCELL_230_1568 ();
 FILLCELL_X32 FILLCELL_230_1600 ();
 FILLCELL_X32 FILLCELL_230_1632 ();
 FILLCELL_X32 FILLCELL_230_1664 ();
 FILLCELL_X32 FILLCELL_230_1696 ();
 FILLCELL_X32 FILLCELL_230_1728 ();
 FILLCELL_X32 FILLCELL_230_1760 ();
 FILLCELL_X32 FILLCELL_230_1792 ();
 FILLCELL_X32 FILLCELL_230_1824 ();
 FILLCELL_X32 FILLCELL_230_1856 ();
 FILLCELL_X8 FILLCELL_230_1888 ();
 FILLCELL_X1 FILLCELL_230_1896 ();
 FILLCELL_X32 FILLCELL_231_0 ();
 FILLCELL_X32 FILLCELL_231_32 ();
 FILLCELL_X32 FILLCELL_231_64 ();
 FILLCELL_X32 FILLCELL_231_96 ();
 FILLCELL_X32 FILLCELL_231_128 ();
 FILLCELL_X32 FILLCELL_231_160 ();
 FILLCELL_X32 FILLCELL_231_192 ();
 FILLCELL_X32 FILLCELL_231_224 ();
 FILLCELL_X32 FILLCELL_231_256 ();
 FILLCELL_X32 FILLCELL_231_288 ();
 FILLCELL_X32 FILLCELL_231_320 ();
 FILLCELL_X32 FILLCELL_231_352 ();
 FILLCELL_X32 FILLCELL_231_384 ();
 FILLCELL_X32 FILLCELL_231_416 ();
 FILLCELL_X32 FILLCELL_231_448 ();
 FILLCELL_X32 FILLCELL_231_480 ();
 FILLCELL_X32 FILLCELL_231_512 ();
 FILLCELL_X32 FILLCELL_231_544 ();
 FILLCELL_X32 FILLCELL_231_576 ();
 FILLCELL_X32 FILLCELL_231_608 ();
 FILLCELL_X32 FILLCELL_231_640 ();
 FILLCELL_X32 FILLCELL_231_672 ();
 FILLCELL_X32 FILLCELL_231_704 ();
 FILLCELL_X32 FILLCELL_231_736 ();
 FILLCELL_X32 FILLCELL_231_768 ();
 FILLCELL_X32 FILLCELL_231_800 ();
 FILLCELL_X32 FILLCELL_231_832 ();
 FILLCELL_X32 FILLCELL_231_864 ();
 FILLCELL_X32 FILLCELL_231_896 ();
 FILLCELL_X32 FILLCELL_231_928 ();
 FILLCELL_X32 FILLCELL_231_960 ();
 FILLCELL_X32 FILLCELL_231_992 ();
 FILLCELL_X32 FILLCELL_231_1024 ();
 FILLCELL_X32 FILLCELL_231_1056 ();
 FILLCELL_X32 FILLCELL_231_1088 ();
 FILLCELL_X32 FILLCELL_231_1120 ();
 FILLCELL_X32 FILLCELL_231_1152 ();
 FILLCELL_X32 FILLCELL_231_1184 ();
 FILLCELL_X32 FILLCELL_231_1216 ();
 FILLCELL_X32 FILLCELL_231_1248 ();
 FILLCELL_X32 FILLCELL_231_1280 ();
 FILLCELL_X32 FILLCELL_231_1312 ();
 FILLCELL_X32 FILLCELL_231_1344 ();
 FILLCELL_X32 FILLCELL_231_1376 ();
 FILLCELL_X32 FILLCELL_231_1408 ();
 FILLCELL_X32 FILLCELL_231_1440 ();
 FILLCELL_X32 FILLCELL_231_1472 ();
 FILLCELL_X32 FILLCELL_231_1504 ();
 FILLCELL_X32 FILLCELL_231_1536 ();
 FILLCELL_X32 FILLCELL_231_1568 ();
 FILLCELL_X32 FILLCELL_231_1600 ();
 FILLCELL_X32 FILLCELL_231_1632 ();
 FILLCELL_X32 FILLCELL_231_1664 ();
 FILLCELL_X32 FILLCELL_231_1696 ();
 FILLCELL_X32 FILLCELL_231_1728 ();
 FILLCELL_X32 FILLCELL_231_1760 ();
 FILLCELL_X32 FILLCELL_231_1792 ();
 FILLCELL_X32 FILLCELL_231_1824 ();
 FILLCELL_X32 FILLCELL_231_1856 ();
 FILLCELL_X8 FILLCELL_231_1888 ();
 FILLCELL_X1 FILLCELL_231_1896 ();
 FILLCELL_X32 FILLCELL_232_0 ();
 FILLCELL_X32 FILLCELL_232_32 ();
 FILLCELL_X32 FILLCELL_232_64 ();
 FILLCELL_X32 FILLCELL_232_96 ();
 FILLCELL_X32 FILLCELL_232_128 ();
 FILLCELL_X32 FILLCELL_232_160 ();
 FILLCELL_X32 FILLCELL_232_192 ();
 FILLCELL_X32 FILLCELL_232_224 ();
 FILLCELL_X32 FILLCELL_232_256 ();
 FILLCELL_X32 FILLCELL_232_288 ();
 FILLCELL_X32 FILLCELL_232_320 ();
 FILLCELL_X32 FILLCELL_232_352 ();
 FILLCELL_X32 FILLCELL_232_384 ();
 FILLCELL_X32 FILLCELL_232_416 ();
 FILLCELL_X32 FILLCELL_232_448 ();
 FILLCELL_X32 FILLCELL_232_480 ();
 FILLCELL_X32 FILLCELL_232_512 ();
 FILLCELL_X32 FILLCELL_232_544 ();
 FILLCELL_X32 FILLCELL_232_576 ();
 FILLCELL_X32 FILLCELL_232_608 ();
 FILLCELL_X32 FILLCELL_232_640 ();
 FILLCELL_X32 FILLCELL_232_672 ();
 FILLCELL_X32 FILLCELL_232_704 ();
 FILLCELL_X32 FILLCELL_232_736 ();
 FILLCELL_X32 FILLCELL_232_768 ();
 FILLCELL_X32 FILLCELL_232_800 ();
 FILLCELL_X32 FILLCELL_232_832 ();
 FILLCELL_X32 FILLCELL_232_864 ();
 FILLCELL_X32 FILLCELL_232_896 ();
 FILLCELL_X32 FILLCELL_232_928 ();
 FILLCELL_X32 FILLCELL_232_960 ();
 FILLCELL_X32 FILLCELL_232_992 ();
 FILLCELL_X32 FILLCELL_232_1024 ();
 FILLCELL_X32 FILLCELL_232_1056 ();
 FILLCELL_X32 FILLCELL_232_1088 ();
 FILLCELL_X32 FILLCELL_232_1120 ();
 FILLCELL_X32 FILLCELL_232_1152 ();
 FILLCELL_X32 FILLCELL_232_1184 ();
 FILLCELL_X32 FILLCELL_232_1216 ();
 FILLCELL_X32 FILLCELL_232_1248 ();
 FILLCELL_X32 FILLCELL_232_1280 ();
 FILLCELL_X32 FILLCELL_232_1312 ();
 FILLCELL_X32 FILLCELL_232_1344 ();
 FILLCELL_X32 FILLCELL_232_1376 ();
 FILLCELL_X32 FILLCELL_232_1408 ();
 FILLCELL_X32 FILLCELL_232_1440 ();
 FILLCELL_X32 FILLCELL_232_1472 ();
 FILLCELL_X32 FILLCELL_232_1504 ();
 FILLCELL_X32 FILLCELL_232_1536 ();
 FILLCELL_X32 FILLCELL_232_1568 ();
 FILLCELL_X32 FILLCELL_232_1600 ();
 FILLCELL_X32 FILLCELL_232_1632 ();
 FILLCELL_X32 FILLCELL_232_1664 ();
 FILLCELL_X32 FILLCELL_232_1696 ();
 FILLCELL_X32 FILLCELL_232_1728 ();
 FILLCELL_X32 FILLCELL_232_1760 ();
 FILLCELL_X32 FILLCELL_232_1792 ();
 FILLCELL_X32 FILLCELL_232_1824 ();
 FILLCELL_X32 FILLCELL_232_1856 ();
 FILLCELL_X8 FILLCELL_232_1888 ();
 FILLCELL_X1 FILLCELL_232_1896 ();
 FILLCELL_X32 FILLCELL_233_0 ();
 FILLCELL_X32 FILLCELL_233_32 ();
 FILLCELL_X32 FILLCELL_233_64 ();
 FILLCELL_X32 FILLCELL_233_96 ();
 FILLCELL_X32 FILLCELL_233_128 ();
 FILLCELL_X32 FILLCELL_233_160 ();
 FILLCELL_X32 FILLCELL_233_192 ();
 FILLCELL_X32 FILLCELL_233_224 ();
 FILLCELL_X32 FILLCELL_233_256 ();
 FILLCELL_X32 FILLCELL_233_288 ();
 FILLCELL_X32 FILLCELL_233_320 ();
 FILLCELL_X32 FILLCELL_233_352 ();
 FILLCELL_X32 FILLCELL_233_384 ();
 FILLCELL_X32 FILLCELL_233_416 ();
 FILLCELL_X32 FILLCELL_233_448 ();
 FILLCELL_X32 FILLCELL_233_480 ();
 FILLCELL_X32 FILLCELL_233_512 ();
 FILLCELL_X32 FILLCELL_233_544 ();
 FILLCELL_X32 FILLCELL_233_576 ();
 FILLCELL_X32 FILLCELL_233_608 ();
 FILLCELL_X32 FILLCELL_233_640 ();
 FILLCELL_X32 FILLCELL_233_672 ();
 FILLCELL_X32 FILLCELL_233_704 ();
 FILLCELL_X32 FILLCELL_233_736 ();
 FILLCELL_X32 FILLCELL_233_768 ();
 FILLCELL_X32 FILLCELL_233_800 ();
 FILLCELL_X32 FILLCELL_233_832 ();
 FILLCELL_X32 FILLCELL_233_864 ();
 FILLCELL_X32 FILLCELL_233_896 ();
 FILLCELL_X32 FILLCELL_233_928 ();
 FILLCELL_X32 FILLCELL_233_960 ();
 FILLCELL_X32 FILLCELL_233_992 ();
 FILLCELL_X32 FILLCELL_233_1024 ();
 FILLCELL_X32 FILLCELL_233_1056 ();
 FILLCELL_X32 FILLCELL_233_1088 ();
 FILLCELL_X32 FILLCELL_233_1120 ();
 FILLCELL_X32 FILLCELL_233_1152 ();
 FILLCELL_X32 FILLCELL_233_1184 ();
 FILLCELL_X32 FILLCELL_233_1216 ();
 FILLCELL_X32 FILLCELL_233_1248 ();
 FILLCELL_X32 FILLCELL_233_1280 ();
 FILLCELL_X32 FILLCELL_233_1312 ();
 FILLCELL_X32 FILLCELL_233_1344 ();
 FILLCELL_X32 FILLCELL_233_1376 ();
 FILLCELL_X32 FILLCELL_233_1408 ();
 FILLCELL_X32 FILLCELL_233_1440 ();
 FILLCELL_X32 FILLCELL_233_1472 ();
 FILLCELL_X32 FILLCELL_233_1504 ();
 FILLCELL_X32 FILLCELL_233_1536 ();
 FILLCELL_X32 FILLCELL_233_1568 ();
 FILLCELL_X32 FILLCELL_233_1600 ();
 FILLCELL_X32 FILLCELL_233_1632 ();
 FILLCELL_X32 FILLCELL_233_1664 ();
 FILLCELL_X32 FILLCELL_233_1696 ();
 FILLCELL_X32 FILLCELL_233_1728 ();
 FILLCELL_X32 FILLCELL_233_1760 ();
 FILLCELL_X32 FILLCELL_233_1792 ();
 FILLCELL_X32 FILLCELL_233_1824 ();
 FILLCELL_X32 FILLCELL_233_1856 ();
 FILLCELL_X8 FILLCELL_233_1888 ();
 FILLCELL_X1 FILLCELL_233_1896 ();
 FILLCELL_X32 FILLCELL_234_0 ();
 FILLCELL_X32 FILLCELL_234_32 ();
 FILLCELL_X32 FILLCELL_234_64 ();
 FILLCELL_X32 FILLCELL_234_96 ();
 FILLCELL_X32 FILLCELL_234_128 ();
 FILLCELL_X32 FILLCELL_234_160 ();
 FILLCELL_X32 FILLCELL_234_192 ();
 FILLCELL_X32 FILLCELL_234_224 ();
 FILLCELL_X32 FILLCELL_234_256 ();
 FILLCELL_X32 FILLCELL_234_288 ();
 FILLCELL_X32 FILLCELL_234_320 ();
 FILLCELL_X32 FILLCELL_234_352 ();
 FILLCELL_X32 FILLCELL_234_384 ();
 FILLCELL_X32 FILLCELL_234_416 ();
 FILLCELL_X32 FILLCELL_234_448 ();
 FILLCELL_X32 FILLCELL_234_480 ();
 FILLCELL_X32 FILLCELL_234_512 ();
 FILLCELL_X32 FILLCELL_234_544 ();
 FILLCELL_X32 FILLCELL_234_576 ();
 FILLCELL_X32 FILLCELL_234_608 ();
 FILLCELL_X32 FILLCELL_234_640 ();
 FILLCELL_X32 FILLCELL_234_672 ();
 FILLCELL_X32 FILLCELL_234_704 ();
 FILLCELL_X32 FILLCELL_234_736 ();
 FILLCELL_X32 FILLCELL_234_768 ();
 FILLCELL_X32 FILLCELL_234_800 ();
 FILLCELL_X32 FILLCELL_234_832 ();
 FILLCELL_X32 FILLCELL_234_864 ();
 FILLCELL_X32 FILLCELL_234_896 ();
 FILLCELL_X32 FILLCELL_234_928 ();
 FILLCELL_X32 FILLCELL_234_960 ();
 FILLCELL_X32 FILLCELL_234_992 ();
 FILLCELL_X32 FILLCELL_234_1024 ();
 FILLCELL_X32 FILLCELL_234_1056 ();
 FILLCELL_X32 FILLCELL_234_1088 ();
 FILLCELL_X32 FILLCELL_234_1120 ();
 FILLCELL_X32 FILLCELL_234_1152 ();
 FILLCELL_X32 FILLCELL_234_1184 ();
 FILLCELL_X32 FILLCELL_234_1216 ();
 FILLCELL_X32 FILLCELL_234_1248 ();
 FILLCELL_X32 FILLCELL_234_1280 ();
 FILLCELL_X32 FILLCELL_234_1312 ();
 FILLCELL_X32 FILLCELL_234_1344 ();
 FILLCELL_X32 FILLCELL_234_1376 ();
 FILLCELL_X32 FILLCELL_234_1408 ();
 FILLCELL_X32 FILLCELL_234_1440 ();
 FILLCELL_X32 FILLCELL_234_1472 ();
 FILLCELL_X32 FILLCELL_234_1504 ();
 FILLCELL_X32 FILLCELL_234_1536 ();
 FILLCELL_X32 FILLCELL_234_1568 ();
 FILLCELL_X32 FILLCELL_234_1600 ();
 FILLCELL_X32 FILLCELL_234_1632 ();
 FILLCELL_X32 FILLCELL_234_1664 ();
 FILLCELL_X32 FILLCELL_234_1696 ();
 FILLCELL_X32 FILLCELL_234_1728 ();
 FILLCELL_X32 FILLCELL_234_1760 ();
 FILLCELL_X32 FILLCELL_234_1792 ();
 FILLCELL_X32 FILLCELL_234_1824 ();
 FILLCELL_X32 FILLCELL_234_1856 ();
 FILLCELL_X8 FILLCELL_234_1888 ();
 FILLCELL_X1 FILLCELL_234_1896 ();
 FILLCELL_X32 FILLCELL_235_0 ();
 FILLCELL_X32 FILLCELL_235_32 ();
 FILLCELL_X32 FILLCELL_235_64 ();
 FILLCELL_X32 FILLCELL_235_96 ();
 FILLCELL_X32 FILLCELL_235_128 ();
 FILLCELL_X32 FILLCELL_235_160 ();
 FILLCELL_X32 FILLCELL_235_192 ();
 FILLCELL_X32 FILLCELL_235_224 ();
 FILLCELL_X32 FILLCELL_235_256 ();
 FILLCELL_X32 FILLCELL_235_288 ();
 FILLCELL_X32 FILLCELL_235_320 ();
 FILLCELL_X32 FILLCELL_235_352 ();
 FILLCELL_X32 FILLCELL_235_384 ();
 FILLCELL_X32 FILLCELL_235_416 ();
 FILLCELL_X32 FILLCELL_235_448 ();
 FILLCELL_X32 FILLCELL_235_480 ();
 FILLCELL_X32 FILLCELL_235_512 ();
 FILLCELL_X32 FILLCELL_235_544 ();
 FILLCELL_X32 FILLCELL_235_576 ();
 FILLCELL_X32 FILLCELL_235_608 ();
 FILLCELL_X32 FILLCELL_235_640 ();
 FILLCELL_X32 FILLCELL_235_672 ();
 FILLCELL_X32 FILLCELL_235_704 ();
 FILLCELL_X32 FILLCELL_235_736 ();
 FILLCELL_X32 FILLCELL_235_768 ();
 FILLCELL_X32 FILLCELL_235_800 ();
 FILLCELL_X32 FILLCELL_235_832 ();
 FILLCELL_X32 FILLCELL_235_864 ();
 FILLCELL_X32 FILLCELL_235_896 ();
 FILLCELL_X32 FILLCELL_235_928 ();
 FILLCELL_X32 FILLCELL_235_960 ();
 FILLCELL_X32 FILLCELL_235_992 ();
 FILLCELL_X32 FILLCELL_235_1024 ();
 FILLCELL_X32 FILLCELL_235_1056 ();
 FILLCELL_X32 FILLCELL_235_1088 ();
 FILLCELL_X32 FILLCELL_235_1120 ();
 FILLCELL_X32 FILLCELL_235_1152 ();
 FILLCELL_X32 FILLCELL_235_1184 ();
 FILLCELL_X32 FILLCELL_235_1216 ();
 FILLCELL_X32 FILLCELL_235_1248 ();
 FILLCELL_X32 FILLCELL_235_1280 ();
 FILLCELL_X32 FILLCELL_235_1312 ();
 FILLCELL_X32 FILLCELL_235_1344 ();
 FILLCELL_X32 FILLCELL_235_1376 ();
 FILLCELL_X32 FILLCELL_235_1408 ();
 FILLCELL_X32 FILLCELL_235_1440 ();
 FILLCELL_X32 FILLCELL_235_1472 ();
 FILLCELL_X32 FILLCELL_235_1504 ();
 FILLCELL_X32 FILLCELL_235_1536 ();
 FILLCELL_X32 FILLCELL_235_1568 ();
 FILLCELL_X32 FILLCELL_235_1600 ();
 FILLCELL_X32 FILLCELL_235_1632 ();
 FILLCELL_X32 FILLCELL_235_1664 ();
 FILLCELL_X32 FILLCELL_235_1696 ();
 FILLCELL_X32 FILLCELL_235_1728 ();
 FILLCELL_X32 FILLCELL_235_1760 ();
 FILLCELL_X32 FILLCELL_235_1792 ();
 FILLCELL_X32 FILLCELL_235_1824 ();
 FILLCELL_X32 FILLCELL_235_1856 ();
 FILLCELL_X8 FILLCELL_235_1888 ();
 FILLCELL_X1 FILLCELL_235_1896 ();
 FILLCELL_X32 FILLCELL_236_0 ();
 FILLCELL_X32 FILLCELL_236_32 ();
 FILLCELL_X32 FILLCELL_236_64 ();
 FILLCELL_X32 FILLCELL_236_96 ();
 FILLCELL_X32 FILLCELL_236_128 ();
 FILLCELL_X32 FILLCELL_236_160 ();
 FILLCELL_X32 FILLCELL_236_192 ();
 FILLCELL_X32 FILLCELL_236_224 ();
 FILLCELL_X32 FILLCELL_236_256 ();
 FILLCELL_X32 FILLCELL_236_288 ();
 FILLCELL_X32 FILLCELL_236_320 ();
 FILLCELL_X32 FILLCELL_236_352 ();
 FILLCELL_X32 FILLCELL_236_384 ();
 FILLCELL_X32 FILLCELL_236_416 ();
 FILLCELL_X32 FILLCELL_236_448 ();
 FILLCELL_X32 FILLCELL_236_480 ();
 FILLCELL_X32 FILLCELL_236_512 ();
 FILLCELL_X32 FILLCELL_236_544 ();
 FILLCELL_X32 FILLCELL_236_576 ();
 FILLCELL_X32 FILLCELL_236_608 ();
 FILLCELL_X32 FILLCELL_236_640 ();
 FILLCELL_X32 FILLCELL_236_672 ();
 FILLCELL_X32 FILLCELL_236_704 ();
 FILLCELL_X32 FILLCELL_236_736 ();
 FILLCELL_X32 FILLCELL_236_768 ();
 FILLCELL_X32 FILLCELL_236_800 ();
 FILLCELL_X32 FILLCELL_236_832 ();
 FILLCELL_X32 FILLCELL_236_864 ();
 FILLCELL_X32 FILLCELL_236_896 ();
 FILLCELL_X32 FILLCELL_236_928 ();
 FILLCELL_X32 FILLCELL_236_960 ();
 FILLCELL_X32 FILLCELL_236_992 ();
 FILLCELL_X32 FILLCELL_236_1024 ();
 FILLCELL_X32 FILLCELL_236_1056 ();
 FILLCELL_X32 FILLCELL_236_1088 ();
 FILLCELL_X32 FILLCELL_236_1120 ();
 FILLCELL_X32 FILLCELL_236_1152 ();
 FILLCELL_X32 FILLCELL_236_1184 ();
 FILLCELL_X32 FILLCELL_236_1216 ();
 FILLCELL_X32 FILLCELL_236_1248 ();
 FILLCELL_X32 FILLCELL_236_1280 ();
 FILLCELL_X32 FILLCELL_236_1312 ();
 FILLCELL_X32 FILLCELL_236_1344 ();
 FILLCELL_X32 FILLCELL_236_1376 ();
 FILLCELL_X32 FILLCELL_236_1408 ();
 FILLCELL_X32 FILLCELL_236_1440 ();
 FILLCELL_X32 FILLCELL_236_1472 ();
 FILLCELL_X32 FILLCELL_236_1504 ();
 FILLCELL_X32 FILLCELL_236_1536 ();
 FILLCELL_X32 FILLCELL_236_1568 ();
 FILLCELL_X32 FILLCELL_236_1600 ();
 FILLCELL_X32 FILLCELL_236_1632 ();
 FILLCELL_X32 FILLCELL_236_1664 ();
 FILLCELL_X32 FILLCELL_236_1696 ();
 FILLCELL_X32 FILLCELL_236_1728 ();
 FILLCELL_X32 FILLCELL_236_1760 ();
 FILLCELL_X32 FILLCELL_236_1792 ();
 FILLCELL_X32 FILLCELL_236_1824 ();
 FILLCELL_X32 FILLCELL_236_1856 ();
 FILLCELL_X8 FILLCELL_236_1888 ();
 FILLCELL_X1 FILLCELL_236_1896 ();
 FILLCELL_X32 FILLCELL_237_0 ();
 FILLCELL_X32 FILLCELL_237_32 ();
 FILLCELL_X32 FILLCELL_237_64 ();
 FILLCELL_X32 FILLCELL_237_96 ();
 FILLCELL_X32 FILLCELL_237_128 ();
 FILLCELL_X32 FILLCELL_237_160 ();
 FILLCELL_X32 FILLCELL_237_192 ();
 FILLCELL_X32 FILLCELL_237_224 ();
 FILLCELL_X32 FILLCELL_237_256 ();
 FILLCELL_X32 FILLCELL_237_288 ();
 FILLCELL_X32 FILLCELL_237_320 ();
 FILLCELL_X32 FILLCELL_237_352 ();
 FILLCELL_X32 FILLCELL_237_384 ();
 FILLCELL_X32 FILLCELL_237_416 ();
 FILLCELL_X32 FILLCELL_237_448 ();
 FILLCELL_X32 FILLCELL_237_480 ();
 FILLCELL_X32 FILLCELL_237_512 ();
 FILLCELL_X32 FILLCELL_237_544 ();
 FILLCELL_X32 FILLCELL_237_576 ();
 FILLCELL_X32 FILLCELL_237_608 ();
 FILLCELL_X32 FILLCELL_237_640 ();
 FILLCELL_X32 FILLCELL_237_672 ();
 FILLCELL_X32 FILLCELL_237_704 ();
 FILLCELL_X32 FILLCELL_237_736 ();
 FILLCELL_X32 FILLCELL_237_768 ();
 FILLCELL_X32 FILLCELL_237_800 ();
 FILLCELL_X32 FILLCELL_237_832 ();
 FILLCELL_X32 FILLCELL_237_864 ();
 FILLCELL_X32 FILLCELL_237_896 ();
 FILLCELL_X32 FILLCELL_237_928 ();
 FILLCELL_X32 FILLCELL_237_960 ();
 FILLCELL_X32 FILLCELL_237_992 ();
 FILLCELL_X32 FILLCELL_237_1024 ();
 FILLCELL_X32 FILLCELL_237_1056 ();
 FILLCELL_X32 FILLCELL_237_1088 ();
 FILLCELL_X32 FILLCELL_237_1120 ();
 FILLCELL_X32 FILLCELL_237_1152 ();
 FILLCELL_X32 FILLCELL_237_1184 ();
 FILLCELL_X32 FILLCELL_237_1216 ();
 FILLCELL_X32 FILLCELL_237_1248 ();
 FILLCELL_X32 FILLCELL_237_1280 ();
 FILLCELL_X32 FILLCELL_237_1312 ();
 FILLCELL_X32 FILLCELL_237_1344 ();
 FILLCELL_X32 FILLCELL_237_1376 ();
 FILLCELL_X32 FILLCELL_237_1408 ();
 FILLCELL_X32 FILLCELL_237_1440 ();
 FILLCELL_X32 FILLCELL_237_1472 ();
 FILLCELL_X32 FILLCELL_237_1504 ();
 FILLCELL_X32 FILLCELL_237_1536 ();
 FILLCELL_X32 FILLCELL_237_1568 ();
 FILLCELL_X32 FILLCELL_237_1600 ();
 FILLCELL_X32 FILLCELL_237_1632 ();
 FILLCELL_X32 FILLCELL_237_1664 ();
 FILLCELL_X32 FILLCELL_237_1696 ();
 FILLCELL_X32 FILLCELL_237_1728 ();
 FILLCELL_X32 FILLCELL_237_1760 ();
 FILLCELL_X32 FILLCELL_237_1792 ();
 FILLCELL_X32 FILLCELL_237_1824 ();
 FILLCELL_X32 FILLCELL_237_1856 ();
 FILLCELL_X8 FILLCELL_237_1888 ();
 FILLCELL_X1 FILLCELL_237_1896 ();
 FILLCELL_X32 FILLCELL_238_0 ();
 FILLCELL_X32 FILLCELL_238_32 ();
 FILLCELL_X32 FILLCELL_238_64 ();
 FILLCELL_X32 FILLCELL_238_96 ();
 FILLCELL_X32 FILLCELL_238_128 ();
 FILLCELL_X32 FILLCELL_238_160 ();
 FILLCELL_X32 FILLCELL_238_192 ();
 FILLCELL_X32 FILLCELL_238_224 ();
 FILLCELL_X32 FILLCELL_238_256 ();
 FILLCELL_X32 FILLCELL_238_288 ();
 FILLCELL_X32 FILLCELL_238_320 ();
 FILLCELL_X32 FILLCELL_238_352 ();
 FILLCELL_X32 FILLCELL_238_384 ();
 FILLCELL_X32 FILLCELL_238_416 ();
 FILLCELL_X32 FILLCELL_238_448 ();
 FILLCELL_X32 FILLCELL_238_480 ();
 FILLCELL_X32 FILLCELL_238_512 ();
 FILLCELL_X32 FILLCELL_238_544 ();
 FILLCELL_X32 FILLCELL_238_576 ();
 FILLCELL_X32 FILLCELL_238_608 ();
 FILLCELL_X32 FILLCELL_238_640 ();
 FILLCELL_X32 FILLCELL_238_672 ();
 FILLCELL_X32 FILLCELL_238_704 ();
 FILLCELL_X32 FILLCELL_238_736 ();
 FILLCELL_X32 FILLCELL_238_768 ();
 FILLCELL_X32 FILLCELL_238_800 ();
 FILLCELL_X32 FILLCELL_238_832 ();
 FILLCELL_X32 FILLCELL_238_864 ();
 FILLCELL_X32 FILLCELL_238_896 ();
 FILLCELL_X32 FILLCELL_238_928 ();
 FILLCELL_X32 FILLCELL_238_960 ();
 FILLCELL_X32 FILLCELL_238_992 ();
 FILLCELL_X32 FILLCELL_238_1024 ();
 FILLCELL_X32 FILLCELL_238_1056 ();
 FILLCELL_X32 FILLCELL_238_1088 ();
 FILLCELL_X32 FILLCELL_238_1120 ();
 FILLCELL_X32 FILLCELL_238_1152 ();
 FILLCELL_X32 FILLCELL_238_1184 ();
 FILLCELL_X32 FILLCELL_238_1216 ();
 FILLCELL_X32 FILLCELL_238_1248 ();
 FILLCELL_X32 FILLCELL_238_1280 ();
 FILLCELL_X32 FILLCELL_238_1312 ();
 FILLCELL_X32 FILLCELL_238_1344 ();
 FILLCELL_X32 FILLCELL_238_1376 ();
 FILLCELL_X32 FILLCELL_238_1408 ();
 FILLCELL_X32 FILLCELL_238_1440 ();
 FILLCELL_X32 FILLCELL_238_1472 ();
 FILLCELL_X32 FILLCELL_238_1504 ();
 FILLCELL_X32 FILLCELL_238_1536 ();
 FILLCELL_X32 FILLCELL_238_1568 ();
 FILLCELL_X32 FILLCELL_238_1600 ();
 FILLCELL_X32 FILLCELL_238_1632 ();
 FILLCELL_X32 FILLCELL_238_1664 ();
 FILLCELL_X32 FILLCELL_238_1696 ();
 FILLCELL_X32 FILLCELL_238_1728 ();
 FILLCELL_X32 FILLCELL_238_1760 ();
 FILLCELL_X32 FILLCELL_238_1792 ();
 FILLCELL_X32 FILLCELL_238_1824 ();
 FILLCELL_X32 FILLCELL_238_1856 ();
 FILLCELL_X8 FILLCELL_238_1888 ();
 FILLCELL_X1 FILLCELL_238_1896 ();
 FILLCELL_X32 FILLCELL_239_0 ();
 FILLCELL_X32 FILLCELL_239_32 ();
 FILLCELL_X32 FILLCELL_239_64 ();
 FILLCELL_X32 FILLCELL_239_96 ();
 FILLCELL_X32 FILLCELL_239_128 ();
 FILLCELL_X32 FILLCELL_239_160 ();
 FILLCELL_X32 FILLCELL_239_192 ();
 FILLCELL_X32 FILLCELL_239_224 ();
 FILLCELL_X32 FILLCELL_239_256 ();
 FILLCELL_X32 FILLCELL_239_288 ();
 FILLCELL_X32 FILLCELL_239_320 ();
 FILLCELL_X32 FILLCELL_239_352 ();
 FILLCELL_X32 FILLCELL_239_384 ();
 FILLCELL_X32 FILLCELL_239_416 ();
 FILLCELL_X32 FILLCELL_239_448 ();
 FILLCELL_X32 FILLCELL_239_480 ();
 FILLCELL_X32 FILLCELL_239_512 ();
 FILLCELL_X32 FILLCELL_239_544 ();
 FILLCELL_X32 FILLCELL_239_576 ();
 FILLCELL_X32 FILLCELL_239_608 ();
 FILLCELL_X32 FILLCELL_239_640 ();
 FILLCELL_X32 FILLCELL_239_672 ();
 FILLCELL_X32 FILLCELL_239_704 ();
 FILLCELL_X32 FILLCELL_239_736 ();
 FILLCELL_X32 FILLCELL_239_768 ();
 FILLCELL_X32 FILLCELL_239_800 ();
 FILLCELL_X32 FILLCELL_239_832 ();
 FILLCELL_X32 FILLCELL_239_864 ();
 FILLCELL_X32 FILLCELL_239_896 ();
 FILLCELL_X32 FILLCELL_239_928 ();
 FILLCELL_X32 FILLCELL_239_960 ();
 FILLCELL_X32 FILLCELL_239_992 ();
 FILLCELL_X32 FILLCELL_239_1024 ();
 FILLCELL_X32 FILLCELL_239_1056 ();
 FILLCELL_X32 FILLCELL_239_1088 ();
 FILLCELL_X32 FILLCELL_239_1120 ();
 FILLCELL_X32 FILLCELL_239_1152 ();
 FILLCELL_X32 FILLCELL_239_1184 ();
 FILLCELL_X32 FILLCELL_239_1216 ();
 FILLCELL_X32 FILLCELL_239_1248 ();
 FILLCELL_X32 FILLCELL_239_1280 ();
 FILLCELL_X32 FILLCELL_239_1312 ();
 FILLCELL_X32 FILLCELL_239_1344 ();
 FILLCELL_X32 FILLCELL_239_1376 ();
 FILLCELL_X32 FILLCELL_239_1408 ();
 FILLCELL_X32 FILLCELL_239_1440 ();
 FILLCELL_X32 FILLCELL_239_1472 ();
 FILLCELL_X32 FILLCELL_239_1504 ();
 FILLCELL_X32 FILLCELL_239_1536 ();
 FILLCELL_X32 FILLCELL_239_1568 ();
 FILLCELL_X32 FILLCELL_239_1600 ();
 FILLCELL_X32 FILLCELL_239_1632 ();
 FILLCELL_X32 FILLCELL_239_1664 ();
 FILLCELL_X32 FILLCELL_239_1696 ();
 FILLCELL_X32 FILLCELL_239_1728 ();
 FILLCELL_X32 FILLCELL_239_1760 ();
 FILLCELL_X32 FILLCELL_239_1792 ();
 FILLCELL_X32 FILLCELL_239_1824 ();
 FILLCELL_X32 FILLCELL_239_1856 ();
 FILLCELL_X8 FILLCELL_239_1888 ();
 FILLCELL_X1 FILLCELL_239_1896 ();
 FILLCELL_X32 FILLCELL_240_0 ();
 FILLCELL_X32 FILLCELL_240_32 ();
 FILLCELL_X32 FILLCELL_240_64 ();
 FILLCELL_X32 FILLCELL_240_96 ();
 FILLCELL_X32 FILLCELL_240_128 ();
 FILLCELL_X32 FILLCELL_240_160 ();
 FILLCELL_X32 FILLCELL_240_192 ();
 FILLCELL_X32 FILLCELL_240_224 ();
 FILLCELL_X32 FILLCELL_240_256 ();
 FILLCELL_X32 FILLCELL_240_288 ();
 FILLCELL_X32 FILLCELL_240_320 ();
 FILLCELL_X32 FILLCELL_240_352 ();
 FILLCELL_X32 FILLCELL_240_384 ();
 FILLCELL_X32 FILLCELL_240_416 ();
 FILLCELL_X32 FILLCELL_240_448 ();
 FILLCELL_X32 FILLCELL_240_480 ();
 FILLCELL_X32 FILLCELL_240_512 ();
 FILLCELL_X32 FILLCELL_240_544 ();
 FILLCELL_X32 FILLCELL_240_576 ();
 FILLCELL_X32 FILLCELL_240_608 ();
 FILLCELL_X32 FILLCELL_240_640 ();
 FILLCELL_X32 FILLCELL_240_672 ();
 FILLCELL_X32 FILLCELL_240_704 ();
 FILLCELL_X32 FILLCELL_240_736 ();
 FILLCELL_X32 FILLCELL_240_768 ();
 FILLCELL_X32 FILLCELL_240_800 ();
 FILLCELL_X32 FILLCELL_240_832 ();
 FILLCELL_X32 FILLCELL_240_864 ();
 FILLCELL_X32 FILLCELL_240_896 ();
 FILLCELL_X32 FILLCELL_240_928 ();
 FILLCELL_X32 FILLCELL_240_960 ();
 FILLCELL_X32 FILLCELL_240_992 ();
 FILLCELL_X32 FILLCELL_240_1024 ();
 FILLCELL_X32 FILLCELL_240_1056 ();
 FILLCELL_X32 FILLCELL_240_1088 ();
 FILLCELL_X32 FILLCELL_240_1120 ();
 FILLCELL_X32 FILLCELL_240_1152 ();
 FILLCELL_X32 FILLCELL_240_1184 ();
 FILLCELL_X32 FILLCELL_240_1216 ();
 FILLCELL_X32 FILLCELL_240_1248 ();
 FILLCELL_X32 FILLCELL_240_1280 ();
 FILLCELL_X32 FILLCELL_240_1312 ();
 FILLCELL_X32 FILLCELL_240_1344 ();
 FILLCELL_X32 FILLCELL_240_1376 ();
 FILLCELL_X32 FILLCELL_240_1408 ();
 FILLCELL_X32 FILLCELL_240_1440 ();
 FILLCELL_X32 FILLCELL_240_1472 ();
 FILLCELL_X32 FILLCELL_240_1504 ();
 FILLCELL_X32 FILLCELL_240_1536 ();
 FILLCELL_X32 FILLCELL_240_1568 ();
 FILLCELL_X32 FILLCELL_240_1600 ();
 FILLCELL_X32 FILLCELL_240_1632 ();
 FILLCELL_X32 FILLCELL_240_1664 ();
 FILLCELL_X32 FILLCELL_240_1696 ();
 FILLCELL_X32 FILLCELL_240_1728 ();
 FILLCELL_X32 FILLCELL_240_1760 ();
 FILLCELL_X32 FILLCELL_240_1792 ();
 FILLCELL_X32 FILLCELL_240_1824 ();
 FILLCELL_X32 FILLCELL_240_1856 ();
 FILLCELL_X8 FILLCELL_240_1888 ();
 FILLCELL_X1 FILLCELL_240_1896 ();
 FILLCELL_X32 FILLCELL_241_0 ();
 FILLCELL_X32 FILLCELL_241_32 ();
 FILLCELL_X32 FILLCELL_241_64 ();
 FILLCELL_X32 FILLCELL_241_96 ();
 FILLCELL_X32 FILLCELL_241_128 ();
 FILLCELL_X32 FILLCELL_241_160 ();
 FILLCELL_X32 FILLCELL_241_192 ();
 FILLCELL_X32 FILLCELL_241_224 ();
 FILLCELL_X32 FILLCELL_241_256 ();
 FILLCELL_X32 FILLCELL_241_288 ();
 FILLCELL_X32 FILLCELL_241_320 ();
 FILLCELL_X32 FILLCELL_241_352 ();
 FILLCELL_X32 FILLCELL_241_384 ();
 FILLCELL_X32 FILLCELL_241_416 ();
 FILLCELL_X32 FILLCELL_241_448 ();
 FILLCELL_X32 FILLCELL_241_480 ();
 FILLCELL_X32 FILLCELL_241_512 ();
 FILLCELL_X32 FILLCELL_241_544 ();
 FILLCELL_X32 FILLCELL_241_576 ();
 FILLCELL_X32 FILLCELL_241_608 ();
 FILLCELL_X32 FILLCELL_241_640 ();
 FILLCELL_X32 FILLCELL_241_672 ();
 FILLCELL_X32 FILLCELL_241_704 ();
 FILLCELL_X32 FILLCELL_241_736 ();
 FILLCELL_X32 FILLCELL_241_768 ();
 FILLCELL_X32 FILLCELL_241_800 ();
 FILLCELL_X32 FILLCELL_241_832 ();
 FILLCELL_X32 FILLCELL_241_864 ();
 FILLCELL_X32 FILLCELL_241_896 ();
 FILLCELL_X32 FILLCELL_241_928 ();
 FILLCELL_X32 FILLCELL_241_960 ();
 FILLCELL_X32 FILLCELL_241_992 ();
 FILLCELL_X32 FILLCELL_241_1024 ();
 FILLCELL_X32 FILLCELL_241_1056 ();
 FILLCELL_X32 FILLCELL_241_1088 ();
 FILLCELL_X32 FILLCELL_241_1120 ();
 FILLCELL_X32 FILLCELL_241_1152 ();
 FILLCELL_X32 FILLCELL_241_1184 ();
 FILLCELL_X32 FILLCELL_241_1216 ();
 FILLCELL_X32 FILLCELL_241_1248 ();
 FILLCELL_X32 FILLCELL_241_1280 ();
 FILLCELL_X32 FILLCELL_241_1312 ();
 FILLCELL_X32 FILLCELL_241_1344 ();
 FILLCELL_X32 FILLCELL_241_1376 ();
 FILLCELL_X32 FILLCELL_241_1408 ();
 FILLCELL_X32 FILLCELL_241_1440 ();
 FILLCELL_X32 FILLCELL_241_1472 ();
 FILLCELL_X32 FILLCELL_241_1504 ();
 FILLCELL_X32 FILLCELL_241_1536 ();
 FILLCELL_X32 FILLCELL_241_1568 ();
 FILLCELL_X32 FILLCELL_241_1600 ();
 FILLCELL_X32 FILLCELL_241_1632 ();
 FILLCELL_X32 FILLCELL_241_1664 ();
 FILLCELL_X32 FILLCELL_241_1696 ();
 FILLCELL_X32 FILLCELL_241_1728 ();
 FILLCELL_X32 FILLCELL_241_1760 ();
 FILLCELL_X32 FILLCELL_241_1792 ();
 FILLCELL_X32 FILLCELL_241_1824 ();
 FILLCELL_X32 FILLCELL_241_1856 ();
 FILLCELL_X8 FILLCELL_241_1888 ();
 FILLCELL_X1 FILLCELL_241_1896 ();
 FILLCELL_X32 FILLCELL_242_0 ();
 FILLCELL_X32 FILLCELL_242_32 ();
 FILLCELL_X32 FILLCELL_242_64 ();
 FILLCELL_X32 FILLCELL_242_96 ();
 FILLCELL_X32 FILLCELL_242_128 ();
 FILLCELL_X32 FILLCELL_242_160 ();
 FILLCELL_X32 FILLCELL_242_192 ();
 FILLCELL_X32 FILLCELL_242_224 ();
 FILLCELL_X32 FILLCELL_242_256 ();
 FILLCELL_X32 FILLCELL_242_288 ();
 FILLCELL_X32 FILLCELL_242_320 ();
 FILLCELL_X32 FILLCELL_242_352 ();
 FILLCELL_X32 FILLCELL_242_384 ();
 FILLCELL_X32 FILLCELL_242_416 ();
 FILLCELL_X32 FILLCELL_242_448 ();
 FILLCELL_X32 FILLCELL_242_480 ();
 FILLCELL_X32 FILLCELL_242_512 ();
 FILLCELL_X32 FILLCELL_242_544 ();
 FILLCELL_X32 FILLCELL_242_576 ();
 FILLCELL_X32 FILLCELL_242_608 ();
 FILLCELL_X32 FILLCELL_242_640 ();
 FILLCELL_X32 FILLCELL_242_672 ();
 FILLCELL_X32 FILLCELL_242_704 ();
 FILLCELL_X32 FILLCELL_242_736 ();
 FILLCELL_X32 FILLCELL_242_768 ();
 FILLCELL_X32 FILLCELL_242_800 ();
 FILLCELL_X32 FILLCELL_242_832 ();
 FILLCELL_X32 FILLCELL_242_864 ();
 FILLCELL_X32 FILLCELL_242_896 ();
 FILLCELL_X32 FILLCELL_242_928 ();
 FILLCELL_X32 FILLCELL_242_960 ();
 FILLCELL_X32 FILLCELL_242_992 ();
 FILLCELL_X32 FILLCELL_242_1024 ();
 FILLCELL_X32 FILLCELL_242_1056 ();
 FILLCELL_X32 FILLCELL_242_1088 ();
 FILLCELL_X32 FILLCELL_242_1120 ();
 FILLCELL_X32 FILLCELL_242_1152 ();
 FILLCELL_X32 FILLCELL_242_1184 ();
 FILLCELL_X32 FILLCELL_242_1216 ();
 FILLCELL_X32 FILLCELL_242_1248 ();
 FILLCELL_X32 FILLCELL_242_1280 ();
 FILLCELL_X32 FILLCELL_242_1312 ();
 FILLCELL_X32 FILLCELL_242_1344 ();
 FILLCELL_X32 FILLCELL_242_1376 ();
 FILLCELL_X32 FILLCELL_242_1408 ();
 FILLCELL_X32 FILLCELL_242_1440 ();
 FILLCELL_X32 FILLCELL_242_1472 ();
 FILLCELL_X32 FILLCELL_242_1504 ();
 FILLCELL_X32 FILLCELL_242_1536 ();
 FILLCELL_X32 FILLCELL_242_1568 ();
 FILLCELL_X32 FILLCELL_242_1600 ();
 FILLCELL_X32 FILLCELL_242_1632 ();
 FILLCELL_X32 FILLCELL_242_1664 ();
 FILLCELL_X32 FILLCELL_242_1696 ();
 FILLCELL_X32 FILLCELL_242_1728 ();
 FILLCELL_X32 FILLCELL_242_1760 ();
 FILLCELL_X32 FILLCELL_242_1792 ();
 FILLCELL_X32 FILLCELL_242_1824 ();
 FILLCELL_X32 FILLCELL_242_1856 ();
 FILLCELL_X8 FILLCELL_242_1888 ();
 FILLCELL_X1 FILLCELL_242_1896 ();
 FILLCELL_X32 FILLCELL_243_0 ();
 FILLCELL_X32 FILLCELL_243_32 ();
 FILLCELL_X32 FILLCELL_243_64 ();
 FILLCELL_X32 FILLCELL_243_96 ();
 FILLCELL_X32 FILLCELL_243_128 ();
 FILLCELL_X32 FILLCELL_243_160 ();
 FILLCELL_X32 FILLCELL_243_192 ();
 FILLCELL_X32 FILLCELL_243_224 ();
 FILLCELL_X32 FILLCELL_243_256 ();
 FILLCELL_X32 FILLCELL_243_288 ();
 FILLCELL_X32 FILLCELL_243_320 ();
 FILLCELL_X32 FILLCELL_243_352 ();
 FILLCELL_X32 FILLCELL_243_384 ();
 FILLCELL_X32 FILLCELL_243_416 ();
 FILLCELL_X32 FILLCELL_243_448 ();
 FILLCELL_X32 FILLCELL_243_480 ();
 FILLCELL_X32 FILLCELL_243_512 ();
 FILLCELL_X32 FILLCELL_243_544 ();
 FILLCELL_X32 FILLCELL_243_576 ();
 FILLCELL_X32 FILLCELL_243_608 ();
 FILLCELL_X32 FILLCELL_243_640 ();
 FILLCELL_X32 FILLCELL_243_672 ();
 FILLCELL_X32 FILLCELL_243_704 ();
 FILLCELL_X32 FILLCELL_243_736 ();
 FILLCELL_X32 FILLCELL_243_768 ();
 FILLCELL_X32 FILLCELL_243_800 ();
 FILLCELL_X32 FILLCELL_243_832 ();
 FILLCELL_X32 FILLCELL_243_864 ();
 FILLCELL_X32 FILLCELL_243_896 ();
 FILLCELL_X32 FILLCELL_243_928 ();
 FILLCELL_X32 FILLCELL_243_960 ();
 FILLCELL_X32 FILLCELL_243_992 ();
 FILLCELL_X32 FILLCELL_243_1024 ();
 FILLCELL_X32 FILLCELL_243_1056 ();
 FILLCELL_X32 FILLCELL_243_1088 ();
 FILLCELL_X32 FILLCELL_243_1120 ();
 FILLCELL_X32 FILLCELL_243_1152 ();
 FILLCELL_X32 FILLCELL_243_1184 ();
 FILLCELL_X32 FILLCELL_243_1216 ();
 FILLCELL_X32 FILLCELL_243_1248 ();
 FILLCELL_X32 FILLCELL_243_1280 ();
 FILLCELL_X32 FILLCELL_243_1312 ();
 FILLCELL_X32 FILLCELL_243_1344 ();
 FILLCELL_X32 FILLCELL_243_1376 ();
 FILLCELL_X32 FILLCELL_243_1408 ();
 FILLCELL_X32 FILLCELL_243_1440 ();
 FILLCELL_X32 FILLCELL_243_1472 ();
 FILLCELL_X32 FILLCELL_243_1504 ();
 FILLCELL_X32 FILLCELL_243_1536 ();
 FILLCELL_X32 FILLCELL_243_1568 ();
 FILLCELL_X32 FILLCELL_243_1600 ();
 FILLCELL_X32 FILLCELL_243_1632 ();
 FILLCELL_X32 FILLCELL_243_1664 ();
 FILLCELL_X32 FILLCELL_243_1696 ();
 FILLCELL_X32 FILLCELL_243_1728 ();
 FILLCELL_X32 FILLCELL_243_1760 ();
 FILLCELL_X32 FILLCELL_243_1792 ();
 FILLCELL_X32 FILLCELL_243_1824 ();
 FILLCELL_X32 FILLCELL_243_1856 ();
 FILLCELL_X8 FILLCELL_243_1888 ();
 FILLCELL_X1 FILLCELL_243_1896 ();
 FILLCELL_X32 FILLCELL_244_0 ();
 FILLCELL_X32 FILLCELL_244_32 ();
 FILLCELL_X32 FILLCELL_244_64 ();
 FILLCELL_X32 FILLCELL_244_96 ();
 FILLCELL_X32 FILLCELL_244_128 ();
 FILLCELL_X32 FILLCELL_244_160 ();
 FILLCELL_X32 FILLCELL_244_192 ();
 FILLCELL_X32 FILLCELL_244_224 ();
 FILLCELL_X32 FILLCELL_244_256 ();
 FILLCELL_X32 FILLCELL_244_288 ();
 FILLCELL_X32 FILLCELL_244_320 ();
 FILLCELL_X32 FILLCELL_244_352 ();
 FILLCELL_X32 FILLCELL_244_384 ();
 FILLCELL_X32 FILLCELL_244_416 ();
 FILLCELL_X32 FILLCELL_244_448 ();
 FILLCELL_X32 FILLCELL_244_480 ();
 FILLCELL_X32 FILLCELL_244_512 ();
 FILLCELL_X32 FILLCELL_244_544 ();
 FILLCELL_X32 FILLCELL_244_576 ();
 FILLCELL_X32 FILLCELL_244_608 ();
 FILLCELL_X32 FILLCELL_244_640 ();
 FILLCELL_X32 FILLCELL_244_672 ();
 FILLCELL_X32 FILLCELL_244_704 ();
 FILLCELL_X32 FILLCELL_244_736 ();
 FILLCELL_X32 FILLCELL_244_768 ();
 FILLCELL_X32 FILLCELL_244_800 ();
 FILLCELL_X32 FILLCELL_244_832 ();
 FILLCELL_X32 FILLCELL_244_864 ();
 FILLCELL_X32 FILLCELL_244_896 ();
 FILLCELL_X32 FILLCELL_244_928 ();
 FILLCELL_X32 FILLCELL_244_960 ();
 FILLCELL_X32 FILLCELL_244_992 ();
 FILLCELL_X32 FILLCELL_244_1024 ();
 FILLCELL_X32 FILLCELL_244_1056 ();
 FILLCELL_X32 FILLCELL_244_1088 ();
 FILLCELL_X32 FILLCELL_244_1120 ();
 FILLCELL_X32 FILLCELL_244_1152 ();
 FILLCELL_X32 FILLCELL_244_1184 ();
 FILLCELL_X32 FILLCELL_244_1216 ();
 FILLCELL_X32 FILLCELL_244_1248 ();
 FILLCELL_X32 FILLCELL_244_1280 ();
 FILLCELL_X32 FILLCELL_244_1312 ();
 FILLCELL_X32 FILLCELL_244_1344 ();
 FILLCELL_X32 FILLCELL_244_1376 ();
 FILLCELL_X32 FILLCELL_244_1408 ();
 FILLCELL_X32 FILLCELL_244_1440 ();
 FILLCELL_X32 FILLCELL_244_1472 ();
 FILLCELL_X32 FILLCELL_244_1504 ();
 FILLCELL_X32 FILLCELL_244_1536 ();
 FILLCELL_X32 FILLCELL_244_1568 ();
 FILLCELL_X32 FILLCELL_244_1600 ();
 FILLCELL_X32 FILLCELL_244_1632 ();
 FILLCELL_X32 FILLCELL_244_1664 ();
 FILLCELL_X32 FILLCELL_244_1696 ();
 FILLCELL_X32 FILLCELL_244_1728 ();
 FILLCELL_X32 FILLCELL_244_1760 ();
 FILLCELL_X32 FILLCELL_244_1792 ();
 FILLCELL_X32 FILLCELL_244_1824 ();
 FILLCELL_X32 FILLCELL_244_1856 ();
 FILLCELL_X8 FILLCELL_244_1888 ();
 FILLCELL_X1 FILLCELL_244_1896 ();
 FILLCELL_X32 FILLCELL_245_0 ();
 FILLCELL_X32 FILLCELL_245_32 ();
 FILLCELL_X32 FILLCELL_245_64 ();
 FILLCELL_X32 FILLCELL_245_96 ();
 FILLCELL_X32 FILLCELL_245_128 ();
 FILLCELL_X32 FILLCELL_245_160 ();
 FILLCELL_X32 FILLCELL_245_192 ();
 FILLCELL_X32 FILLCELL_245_224 ();
 FILLCELL_X32 FILLCELL_245_256 ();
 FILLCELL_X32 FILLCELL_245_288 ();
 FILLCELL_X32 FILLCELL_245_320 ();
 FILLCELL_X32 FILLCELL_245_352 ();
 FILLCELL_X32 FILLCELL_245_384 ();
 FILLCELL_X32 FILLCELL_245_416 ();
 FILLCELL_X32 FILLCELL_245_448 ();
 FILLCELL_X32 FILLCELL_245_480 ();
 FILLCELL_X32 FILLCELL_245_512 ();
 FILLCELL_X32 FILLCELL_245_544 ();
 FILLCELL_X32 FILLCELL_245_576 ();
 FILLCELL_X32 FILLCELL_245_608 ();
 FILLCELL_X32 FILLCELL_245_640 ();
 FILLCELL_X32 FILLCELL_245_672 ();
 FILLCELL_X32 FILLCELL_245_704 ();
 FILLCELL_X32 FILLCELL_245_736 ();
 FILLCELL_X32 FILLCELL_245_768 ();
 FILLCELL_X32 FILLCELL_245_800 ();
 FILLCELL_X32 FILLCELL_245_832 ();
 FILLCELL_X32 FILLCELL_245_864 ();
 FILLCELL_X32 FILLCELL_245_896 ();
 FILLCELL_X32 FILLCELL_245_928 ();
 FILLCELL_X32 FILLCELL_245_960 ();
 FILLCELL_X32 FILLCELL_245_992 ();
 FILLCELL_X32 FILLCELL_245_1024 ();
 FILLCELL_X32 FILLCELL_245_1056 ();
 FILLCELL_X32 FILLCELL_245_1088 ();
 FILLCELL_X32 FILLCELL_245_1120 ();
 FILLCELL_X32 FILLCELL_245_1152 ();
 FILLCELL_X32 FILLCELL_245_1184 ();
 FILLCELL_X32 FILLCELL_245_1216 ();
 FILLCELL_X32 FILLCELL_245_1248 ();
 FILLCELL_X32 FILLCELL_245_1280 ();
 FILLCELL_X32 FILLCELL_245_1312 ();
 FILLCELL_X32 FILLCELL_245_1344 ();
 FILLCELL_X32 FILLCELL_245_1376 ();
 FILLCELL_X32 FILLCELL_245_1408 ();
 FILLCELL_X32 FILLCELL_245_1440 ();
 FILLCELL_X32 FILLCELL_245_1472 ();
 FILLCELL_X32 FILLCELL_245_1504 ();
 FILLCELL_X32 FILLCELL_245_1536 ();
 FILLCELL_X32 FILLCELL_245_1568 ();
 FILLCELL_X32 FILLCELL_245_1600 ();
 FILLCELL_X32 FILLCELL_245_1632 ();
 FILLCELL_X32 FILLCELL_245_1664 ();
 FILLCELL_X32 FILLCELL_245_1696 ();
 FILLCELL_X32 FILLCELL_245_1728 ();
 FILLCELL_X32 FILLCELL_245_1760 ();
 FILLCELL_X32 FILLCELL_245_1792 ();
 FILLCELL_X32 FILLCELL_245_1824 ();
 FILLCELL_X32 FILLCELL_245_1856 ();
 FILLCELL_X8 FILLCELL_245_1888 ();
 FILLCELL_X1 FILLCELL_245_1896 ();
 FILLCELL_X32 FILLCELL_246_0 ();
 FILLCELL_X32 FILLCELL_246_32 ();
 FILLCELL_X32 FILLCELL_246_64 ();
 FILLCELL_X32 FILLCELL_246_96 ();
 FILLCELL_X32 FILLCELL_246_128 ();
 FILLCELL_X32 FILLCELL_246_160 ();
 FILLCELL_X32 FILLCELL_246_192 ();
 FILLCELL_X32 FILLCELL_246_224 ();
 FILLCELL_X32 FILLCELL_246_256 ();
 FILLCELL_X32 FILLCELL_246_288 ();
 FILLCELL_X32 FILLCELL_246_320 ();
 FILLCELL_X32 FILLCELL_246_352 ();
 FILLCELL_X32 FILLCELL_246_384 ();
 FILLCELL_X32 FILLCELL_246_416 ();
 FILLCELL_X32 FILLCELL_246_448 ();
 FILLCELL_X32 FILLCELL_246_480 ();
 FILLCELL_X32 FILLCELL_246_512 ();
 FILLCELL_X32 FILLCELL_246_544 ();
 FILLCELL_X32 FILLCELL_246_576 ();
 FILLCELL_X32 FILLCELL_246_608 ();
 FILLCELL_X32 FILLCELL_246_640 ();
 FILLCELL_X32 FILLCELL_246_672 ();
 FILLCELL_X32 FILLCELL_246_704 ();
 FILLCELL_X32 FILLCELL_246_736 ();
 FILLCELL_X32 FILLCELL_246_768 ();
 FILLCELL_X32 FILLCELL_246_800 ();
 FILLCELL_X32 FILLCELL_246_832 ();
 FILLCELL_X32 FILLCELL_246_864 ();
 FILLCELL_X32 FILLCELL_246_896 ();
 FILLCELL_X32 FILLCELL_246_928 ();
 FILLCELL_X32 FILLCELL_246_960 ();
 FILLCELL_X32 FILLCELL_246_992 ();
 FILLCELL_X32 FILLCELL_246_1024 ();
 FILLCELL_X32 FILLCELL_246_1056 ();
 FILLCELL_X32 FILLCELL_246_1088 ();
 FILLCELL_X32 FILLCELL_246_1120 ();
 FILLCELL_X32 FILLCELL_246_1152 ();
 FILLCELL_X32 FILLCELL_246_1184 ();
 FILLCELL_X32 FILLCELL_246_1216 ();
 FILLCELL_X32 FILLCELL_246_1248 ();
 FILLCELL_X32 FILLCELL_246_1280 ();
 FILLCELL_X32 FILLCELL_246_1312 ();
 FILLCELL_X32 FILLCELL_246_1344 ();
 FILLCELL_X32 FILLCELL_246_1376 ();
 FILLCELL_X32 FILLCELL_246_1408 ();
 FILLCELL_X32 FILLCELL_246_1440 ();
 FILLCELL_X32 FILLCELL_246_1472 ();
 FILLCELL_X32 FILLCELL_246_1504 ();
 FILLCELL_X32 FILLCELL_246_1536 ();
 FILLCELL_X32 FILLCELL_246_1568 ();
 FILLCELL_X32 FILLCELL_246_1600 ();
 FILLCELL_X32 FILLCELL_246_1632 ();
 FILLCELL_X32 FILLCELL_246_1664 ();
 FILLCELL_X32 FILLCELL_246_1696 ();
 FILLCELL_X32 FILLCELL_246_1728 ();
 FILLCELL_X32 FILLCELL_246_1760 ();
 FILLCELL_X32 FILLCELL_246_1792 ();
 FILLCELL_X32 FILLCELL_246_1824 ();
 FILLCELL_X32 FILLCELL_246_1856 ();
 FILLCELL_X8 FILLCELL_246_1888 ();
 FILLCELL_X1 FILLCELL_246_1896 ();
 FILLCELL_X32 FILLCELL_247_0 ();
 FILLCELL_X32 FILLCELL_247_32 ();
 FILLCELL_X32 FILLCELL_247_64 ();
 FILLCELL_X32 FILLCELL_247_96 ();
 FILLCELL_X32 FILLCELL_247_128 ();
 FILLCELL_X32 FILLCELL_247_160 ();
 FILLCELL_X32 FILLCELL_247_192 ();
 FILLCELL_X32 FILLCELL_247_224 ();
 FILLCELL_X32 FILLCELL_247_256 ();
 FILLCELL_X32 FILLCELL_247_288 ();
 FILLCELL_X32 FILLCELL_247_320 ();
 FILLCELL_X32 FILLCELL_247_352 ();
 FILLCELL_X32 FILLCELL_247_384 ();
 FILLCELL_X32 FILLCELL_247_416 ();
 FILLCELL_X32 FILLCELL_247_448 ();
 FILLCELL_X32 FILLCELL_247_480 ();
 FILLCELL_X32 FILLCELL_247_512 ();
 FILLCELL_X32 FILLCELL_247_544 ();
 FILLCELL_X32 FILLCELL_247_576 ();
 FILLCELL_X32 FILLCELL_247_608 ();
 FILLCELL_X32 FILLCELL_247_640 ();
 FILLCELL_X32 FILLCELL_247_672 ();
 FILLCELL_X32 FILLCELL_247_704 ();
 FILLCELL_X32 FILLCELL_247_736 ();
 FILLCELL_X32 FILLCELL_247_768 ();
 FILLCELL_X32 FILLCELL_247_800 ();
 FILLCELL_X32 FILLCELL_247_832 ();
 FILLCELL_X32 FILLCELL_247_864 ();
 FILLCELL_X32 FILLCELL_247_896 ();
 FILLCELL_X32 FILLCELL_247_928 ();
 FILLCELL_X32 FILLCELL_247_960 ();
 FILLCELL_X32 FILLCELL_247_992 ();
 FILLCELL_X32 FILLCELL_247_1024 ();
 FILLCELL_X32 FILLCELL_247_1056 ();
 FILLCELL_X32 FILLCELL_247_1088 ();
 FILLCELL_X32 FILLCELL_247_1120 ();
 FILLCELL_X32 FILLCELL_247_1152 ();
 FILLCELL_X32 FILLCELL_247_1184 ();
 FILLCELL_X32 FILLCELL_247_1216 ();
 FILLCELL_X32 FILLCELL_247_1248 ();
 FILLCELL_X32 FILLCELL_247_1280 ();
 FILLCELL_X32 FILLCELL_247_1312 ();
 FILLCELL_X32 FILLCELL_247_1344 ();
 FILLCELL_X32 FILLCELL_247_1376 ();
 FILLCELL_X32 FILLCELL_247_1408 ();
 FILLCELL_X32 FILLCELL_247_1440 ();
 FILLCELL_X32 FILLCELL_247_1472 ();
 FILLCELL_X32 FILLCELL_247_1504 ();
 FILLCELL_X32 FILLCELL_247_1536 ();
 FILLCELL_X32 FILLCELL_247_1568 ();
 FILLCELL_X32 FILLCELL_247_1600 ();
 FILLCELL_X32 FILLCELL_247_1632 ();
 FILLCELL_X32 FILLCELL_247_1664 ();
 FILLCELL_X32 FILLCELL_247_1696 ();
 FILLCELL_X32 FILLCELL_247_1728 ();
 FILLCELL_X32 FILLCELL_247_1760 ();
 FILLCELL_X32 FILLCELL_247_1792 ();
 FILLCELL_X32 FILLCELL_247_1824 ();
 FILLCELL_X32 FILLCELL_247_1856 ();
 FILLCELL_X8 FILLCELL_247_1888 ();
 FILLCELL_X1 FILLCELL_247_1896 ();
 FILLCELL_X32 FILLCELL_248_0 ();
 FILLCELL_X32 FILLCELL_248_32 ();
 FILLCELL_X32 FILLCELL_248_64 ();
 FILLCELL_X32 FILLCELL_248_96 ();
 FILLCELL_X32 FILLCELL_248_128 ();
 FILLCELL_X32 FILLCELL_248_160 ();
 FILLCELL_X32 FILLCELL_248_192 ();
 FILLCELL_X32 FILLCELL_248_224 ();
 FILLCELL_X32 FILLCELL_248_256 ();
 FILLCELL_X32 FILLCELL_248_288 ();
 FILLCELL_X32 FILLCELL_248_320 ();
 FILLCELL_X32 FILLCELL_248_352 ();
 FILLCELL_X32 FILLCELL_248_384 ();
 FILLCELL_X32 FILLCELL_248_416 ();
 FILLCELL_X32 FILLCELL_248_448 ();
 FILLCELL_X32 FILLCELL_248_480 ();
 FILLCELL_X32 FILLCELL_248_512 ();
 FILLCELL_X32 FILLCELL_248_544 ();
 FILLCELL_X32 FILLCELL_248_576 ();
 FILLCELL_X32 FILLCELL_248_608 ();
 FILLCELL_X32 FILLCELL_248_640 ();
 FILLCELL_X32 FILLCELL_248_672 ();
 FILLCELL_X32 FILLCELL_248_704 ();
 FILLCELL_X32 FILLCELL_248_736 ();
 FILLCELL_X32 FILLCELL_248_768 ();
 FILLCELL_X32 FILLCELL_248_800 ();
 FILLCELL_X32 FILLCELL_248_832 ();
 FILLCELL_X32 FILLCELL_248_864 ();
 FILLCELL_X32 FILLCELL_248_896 ();
 FILLCELL_X32 FILLCELL_248_928 ();
 FILLCELL_X32 FILLCELL_248_960 ();
 FILLCELL_X32 FILLCELL_248_992 ();
 FILLCELL_X32 FILLCELL_248_1024 ();
 FILLCELL_X32 FILLCELL_248_1056 ();
 FILLCELL_X32 FILLCELL_248_1088 ();
 FILLCELL_X32 FILLCELL_248_1120 ();
 FILLCELL_X32 FILLCELL_248_1152 ();
 FILLCELL_X32 FILLCELL_248_1184 ();
 FILLCELL_X32 FILLCELL_248_1216 ();
 FILLCELL_X32 FILLCELL_248_1248 ();
 FILLCELL_X32 FILLCELL_248_1280 ();
 FILLCELL_X32 FILLCELL_248_1312 ();
 FILLCELL_X32 FILLCELL_248_1344 ();
 FILLCELL_X32 FILLCELL_248_1376 ();
 FILLCELL_X32 FILLCELL_248_1408 ();
 FILLCELL_X32 FILLCELL_248_1440 ();
 FILLCELL_X32 FILLCELL_248_1472 ();
 FILLCELL_X32 FILLCELL_248_1504 ();
 FILLCELL_X32 FILLCELL_248_1536 ();
 FILLCELL_X32 FILLCELL_248_1568 ();
 FILLCELL_X32 FILLCELL_248_1600 ();
 FILLCELL_X32 FILLCELL_248_1632 ();
 FILLCELL_X32 FILLCELL_248_1664 ();
 FILLCELL_X32 FILLCELL_248_1696 ();
 FILLCELL_X32 FILLCELL_248_1728 ();
 FILLCELL_X32 FILLCELL_248_1760 ();
 FILLCELL_X32 FILLCELL_248_1792 ();
 FILLCELL_X32 FILLCELL_248_1824 ();
 FILLCELL_X32 FILLCELL_248_1856 ();
 FILLCELL_X8 FILLCELL_248_1888 ();
 FILLCELL_X1 FILLCELL_248_1896 ();
 FILLCELL_X32 FILLCELL_249_0 ();
 FILLCELL_X32 FILLCELL_249_32 ();
 FILLCELL_X32 FILLCELL_249_64 ();
 FILLCELL_X32 FILLCELL_249_96 ();
 FILLCELL_X32 FILLCELL_249_128 ();
 FILLCELL_X32 FILLCELL_249_160 ();
 FILLCELL_X32 FILLCELL_249_192 ();
 FILLCELL_X32 FILLCELL_249_224 ();
 FILLCELL_X32 FILLCELL_249_256 ();
 FILLCELL_X32 FILLCELL_249_288 ();
 FILLCELL_X32 FILLCELL_249_320 ();
 FILLCELL_X32 FILLCELL_249_352 ();
 FILLCELL_X32 FILLCELL_249_384 ();
 FILLCELL_X32 FILLCELL_249_416 ();
 FILLCELL_X32 FILLCELL_249_448 ();
 FILLCELL_X32 FILLCELL_249_480 ();
 FILLCELL_X32 FILLCELL_249_512 ();
 FILLCELL_X32 FILLCELL_249_544 ();
 FILLCELL_X32 FILLCELL_249_576 ();
 FILLCELL_X32 FILLCELL_249_608 ();
 FILLCELL_X32 FILLCELL_249_640 ();
 FILLCELL_X32 FILLCELL_249_672 ();
 FILLCELL_X32 FILLCELL_249_704 ();
 FILLCELL_X32 FILLCELL_249_736 ();
 FILLCELL_X32 FILLCELL_249_768 ();
 FILLCELL_X32 FILLCELL_249_800 ();
 FILLCELL_X32 FILLCELL_249_832 ();
 FILLCELL_X32 FILLCELL_249_864 ();
 FILLCELL_X32 FILLCELL_249_896 ();
 FILLCELL_X32 FILLCELL_249_928 ();
 FILLCELL_X32 FILLCELL_249_960 ();
 FILLCELL_X32 FILLCELL_249_992 ();
 FILLCELL_X32 FILLCELL_249_1024 ();
 FILLCELL_X32 FILLCELL_249_1056 ();
 FILLCELL_X32 FILLCELL_249_1088 ();
 FILLCELL_X32 FILLCELL_249_1120 ();
 FILLCELL_X32 FILLCELL_249_1152 ();
 FILLCELL_X32 FILLCELL_249_1184 ();
 FILLCELL_X32 FILLCELL_249_1216 ();
 FILLCELL_X32 FILLCELL_249_1248 ();
 FILLCELL_X32 FILLCELL_249_1280 ();
 FILLCELL_X32 FILLCELL_249_1312 ();
 FILLCELL_X32 FILLCELL_249_1344 ();
 FILLCELL_X32 FILLCELL_249_1376 ();
 FILLCELL_X32 FILLCELL_249_1408 ();
 FILLCELL_X32 FILLCELL_249_1440 ();
 FILLCELL_X32 FILLCELL_249_1472 ();
 FILLCELL_X32 FILLCELL_249_1504 ();
 FILLCELL_X32 FILLCELL_249_1536 ();
 FILLCELL_X32 FILLCELL_249_1568 ();
 FILLCELL_X32 FILLCELL_249_1600 ();
 FILLCELL_X32 FILLCELL_249_1632 ();
 FILLCELL_X32 FILLCELL_249_1664 ();
 FILLCELL_X32 FILLCELL_249_1696 ();
 FILLCELL_X32 FILLCELL_249_1728 ();
 FILLCELL_X32 FILLCELL_249_1760 ();
 FILLCELL_X32 FILLCELL_249_1792 ();
 FILLCELL_X32 FILLCELL_249_1824 ();
 FILLCELL_X32 FILLCELL_249_1856 ();
 FILLCELL_X8 FILLCELL_249_1888 ();
 FILLCELL_X1 FILLCELL_249_1896 ();
 FILLCELL_X32 FILLCELL_250_0 ();
 FILLCELL_X32 FILLCELL_250_32 ();
 FILLCELL_X32 FILLCELL_250_64 ();
 FILLCELL_X32 FILLCELL_250_96 ();
 FILLCELL_X32 FILLCELL_250_128 ();
 FILLCELL_X32 FILLCELL_250_160 ();
 FILLCELL_X32 FILLCELL_250_192 ();
 FILLCELL_X32 FILLCELL_250_224 ();
 FILLCELL_X32 FILLCELL_250_256 ();
 FILLCELL_X32 FILLCELL_250_288 ();
 FILLCELL_X32 FILLCELL_250_320 ();
 FILLCELL_X32 FILLCELL_250_352 ();
 FILLCELL_X32 FILLCELL_250_384 ();
 FILLCELL_X32 FILLCELL_250_416 ();
 FILLCELL_X32 FILLCELL_250_448 ();
 FILLCELL_X32 FILLCELL_250_480 ();
 FILLCELL_X32 FILLCELL_250_512 ();
 FILLCELL_X32 FILLCELL_250_544 ();
 FILLCELL_X32 FILLCELL_250_576 ();
 FILLCELL_X32 FILLCELL_250_608 ();
 FILLCELL_X32 FILLCELL_250_640 ();
 FILLCELL_X32 FILLCELL_250_672 ();
 FILLCELL_X32 FILLCELL_250_704 ();
 FILLCELL_X32 FILLCELL_250_736 ();
 FILLCELL_X32 FILLCELL_250_768 ();
 FILLCELL_X32 FILLCELL_250_800 ();
 FILLCELL_X32 FILLCELL_250_832 ();
 FILLCELL_X32 FILLCELL_250_864 ();
 FILLCELL_X32 FILLCELL_250_896 ();
 FILLCELL_X32 FILLCELL_250_928 ();
 FILLCELL_X32 FILLCELL_250_960 ();
 FILLCELL_X32 FILLCELL_250_992 ();
 FILLCELL_X32 FILLCELL_250_1024 ();
 FILLCELL_X32 FILLCELL_250_1056 ();
 FILLCELL_X32 FILLCELL_250_1088 ();
 FILLCELL_X32 FILLCELL_250_1120 ();
 FILLCELL_X32 FILLCELL_250_1152 ();
 FILLCELL_X32 FILLCELL_250_1184 ();
 FILLCELL_X32 FILLCELL_250_1216 ();
 FILLCELL_X32 FILLCELL_250_1248 ();
 FILLCELL_X32 FILLCELL_250_1280 ();
 FILLCELL_X32 FILLCELL_250_1312 ();
 FILLCELL_X32 FILLCELL_250_1344 ();
 FILLCELL_X32 FILLCELL_250_1376 ();
 FILLCELL_X32 FILLCELL_250_1408 ();
 FILLCELL_X32 FILLCELL_250_1440 ();
 FILLCELL_X32 FILLCELL_250_1472 ();
 FILLCELL_X32 FILLCELL_250_1504 ();
 FILLCELL_X32 FILLCELL_250_1536 ();
 FILLCELL_X32 FILLCELL_250_1568 ();
 FILLCELL_X32 FILLCELL_250_1600 ();
 FILLCELL_X32 FILLCELL_250_1632 ();
 FILLCELL_X32 FILLCELL_250_1664 ();
 FILLCELL_X32 FILLCELL_250_1696 ();
 FILLCELL_X32 FILLCELL_250_1728 ();
 FILLCELL_X32 FILLCELL_250_1760 ();
 FILLCELL_X32 FILLCELL_250_1792 ();
 FILLCELL_X32 FILLCELL_250_1824 ();
 FILLCELL_X32 FILLCELL_250_1856 ();
 FILLCELL_X8 FILLCELL_250_1888 ();
 FILLCELL_X1 FILLCELL_250_1896 ();
 FILLCELL_X32 FILLCELL_251_0 ();
 FILLCELL_X32 FILLCELL_251_32 ();
 FILLCELL_X32 FILLCELL_251_64 ();
 FILLCELL_X32 FILLCELL_251_96 ();
 FILLCELL_X32 FILLCELL_251_128 ();
 FILLCELL_X32 FILLCELL_251_160 ();
 FILLCELL_X32 FILLCELL_251_192 ();
 FILLCELL_X32 FILLCELL_251_224 ();
 FILLCELL_X32 FILLCELL_251_256 ();
 FILLCELL_X32 FILLCELL_251_288 ();
 FILLCELL_X32 FILLCELL_251_320 ();
 FILLCELL_X32 FILLCELL_251_352 ();
 FILLCELL_X32 FILLCELL_251_384 ();
 FILLCELL_X32 FILLCELL_251_416 ();
 FILLCELL_X32 FILLCELL_251_448 ();
 FILLCELL_X32 FILLCELL_251_480 ();
 FILLCELL_X32 FILLCELL_251_512 ();
 FILLCELL_X32 FILLCELL_251_544 ();
 FILLCELL_X32 FILLCELL_251_576 ();
 FILLCELL_X32 FILLCELL_251_608 ();
 FILLCELL_X32 FILLCELL_251_640 ();
 FILLCELL_X32 FILLCELL_251_672 ();
 FILLCELL_X32 FILLCELL_251_704 ();
 FILLCELL_X32 FILLCELL_251_736 ();
 FILLCELL_X32 FILLCELL_251_768 ();
 FILLCELL_X32 FILLCELL_251_800 ();
 FILLCELL_X32 FILLCELL_251_832 ();
 FILLCELL_X32 FILLCELL_251_864 ();
 FILLCELL_X32 FILLCELL_251_896 ();
 FILLCELL_X32 FILLCELL_251_928 ();
 FILLCELL_X32 FILLCELL_251_960 ();
 FILLCELL_X32 FILLCELL_251_992 ();
 FILLCELL_X32 FILLCELL_251_1024 ();
 FILLCELL_X32 FILLCELL_251_1056 ();
 FILLCELL_X32 FILLCELL_251_1088 ();
 FILLCELL_X32 FILLCELL_251_1120 ();
 FILLCELL_X32 FILLCELL_251_1152 ();
 FILLCELL_X32 FILLCELL_251_1184 ();
 FILLCELL_X32 FILLCELL_251_1216 ();
 FILLCELL_X32 FILLCELL_251_1248 ();
 FILLCELL_X32 FILLCELL_251_1280 ();
 FILLCELL_X32 FILLCELL_251_1312 ();
 FILLCELL_X32 FILLCELL_251_1344 ();
 FILLCELL_X32 FILLCELL_251_1376 ();
 FILLCELL_X32 FILLCELL_251_1408 ();
 FILLCELL_X32 FILLCELL_251_1440 ();
 FILLCELL_X32 FILLCELL_251_1472 ();
 FILLCELL_X32 FILLCELL_251_1504 ();
 FILLCELL_X32 FILLCELL_251_1536 ();
 FILLCELL_X32 FILLCELL_251_1568 ();
 FILLCELL_X32 FILLCELL_251_1600 ();
 FILLCELL_X32 FILLCELL_251_1632 ();
 FILLCELL_X32 FILLCELL_251_1664 ();
 FILLCELL_X32 FILLCELL_251_1696 ();
 FILLCELL_X32 FILLCELL_251_1728 ();
 FILLCELL_X32 FILLCELL_251_1760 ();
 FILLCELL_X32 FILLCELL_251_1792 ();
 FILLCELL_X32 FILLCELL_251_1824 ();
 FILLCELL_X32 FILLCELL_251_1856 ();
 FILLCELL_X8 FILLCELL_251_1888 ();
 FILLCELL_X1 FILLCELL_251_1896 ();
 FILLCELL_X32 FILLCELL_252_0 ();
 FILLCELL_X32 FILLCELL_252_32 ();
 FILLCELL_X32 FILLCELL_252_64 ();
 FILLCELL_X32 FILLCELL_252_96 ();
 FILLCELL_X32 FILLCELL_252_128 ();
 FILLCELL_X32 FILLCELL_252_160 ();
 FILLCELL_X32 FILLCELL_252_192 ();
 FILLCELL_X32 FILLCELL_252_224 ();
 FILLCELL_X32 FILLCELL_252_256 ();
 FILLCELL_X32 FILLCELL_252_288 ();
 FILLCELL_X32 FILLCELL_252_320 ();
 FILLCELL_X32 FILLCELL_252_352 ();
 FILLCELL_X32 FILLCELL_252_384 ();
 FILLCELL_X32 FILLCELL_252_416 ();
 FILLCELL_X32 FILLCELL_252_448 ();
 FILLCELL_X32 FILLCELL_252_480 ();
 FILLCELL_X32 FILLCELL_252_512 ();
 FILLCELL_X32 FILLCELL_252_544 ();
 FILLCELL_X32 FILLCELL_252_576 ();
 FILLCELL_X32 FILLCELL_252_608 ();
 FILLCELL_X32 FILLCELL_252_640 ();
 FILLCELL_X32 FILLCELL_252_672 ();
 FILLCELL_X32 FILLCELL_252_704 ();
 FILLCELL_X32 FILLCELL_252_736 ();
 FILLCELL_X32 FILLCELL_252_768 ();
 FILLCELL_X32 FILLCELL_252_800 ();
 FILLCELL_X32 FILLCELL_252_832 ();
 FILLCELL_X32 FILLCELL_252_864 ();
 FILLCELL_X32 FILLCELL_252_896 ();
 FILLCELL_X32 FILLCELL_252_928 ();
 FILLCELL_X32 FILLCELL_252_960 ();
 FILLCELL_X32 FILLCELL_252_992 ();
 FILLCELL_X32 FILLCELL_252_1024 ();
 FILLCELL_X32 FILLCELL_252_1056 ();
 FILLCELL_X32 FILLCELL_252_1088 ();
 FILLCELL_X32 FILLCELL_252_1120 ();
 FILLCELL_X32 FILLCELL_252_1152 ();
 FILLCELL_X32 FILLCELL_252_1184 ();
 FILLCELL_X32 FILLCELL_252_1216 ();
 FILLCELL_X32 FILLCELL_252_1248 ();
 FILLCELL_X32 FILLCELL_252_1280 ();
 FILLCELL_X32 FILLCELL_252_1312 ();
 FILLCELL_X32 FILLCELL_252_1344 ();
 FILLCELL_X32 FILLCELL_252_1376 ();
 FILLCELL_X32 FILLCELL_252_1408 ();
 FILLCELL_X32 FILLCELL_252_1440 ();
 FILLCELL_X32 FILLCELL_252_1472 ();
 FILLCELL_X32 FILLCELL_252_1504 ();
 FILLCELL_X32 FILLCELL_252_1536 ();
 FILLCELL_X32 FILLCELL_252_1568 ();
 FILLCELL_X32 FILLCELL_252_1600 ();
 FILLCELL_X32 FILLCELL_252_1632 ();
 FILLCELL_X32 FILLCELL_252_1664 ();
 FILLCELL_X32 FILLCELL_252_1696 ();
 FILLCELL_X32 FILLCELL_252_1728 ();
 FILLCELL_X32 FILLCELL_252_1760 ();
 FILLCELL_X32 FILLCELL_252_1792 ();
 FILLCELL_X32 FILLCELL_252_1824 ();
 FILLCELL_X32 FILLCELL_252_1856 ();
 FILLCELL_X8 FILLCELL_252_1888 ();
 FILLCELL_X1 FILLCELL_252_1896 ();
 FILLCELL_X32 FILLCELL_253_0 ();
 FILLCELL_X32 FILLCELL_253_32 ();
 FILLCELL_X32 FILLCELL_253_64 ();
 FILLCELL_X32 FILLCELL_253_96 ();
 FILLCELL_X32 FILLCELL_253_128 ();
 FILLCELL_X32 FILLCELL_253_160 ();
 FILLCELL_X32 FILLCELL_253_192 ();
 FILLCELL_X32 FILLCELL_253_224 ();
 FILLCELL_X32 FILLCELL_253_256 ();
 FILLCELL_X32 FILLCELL_253_288 ();
 FILLCELL_X32 FILLCELL_253_320 ();
 FILLCELL_X32 FILLCELL_253_352 ();
 FILLCELL_X32 FILLCELL_253_384 ();
 FILLCELL_X32 FILLCELL_253_416 ();
 FILLCELL_X32 FILLCELL_253_448 ();
 FILLCELL_X32 FILLCELL_253_480 ();
 FILLCELL_X32 FILLCELL_253_512 ();
 FILLCELL_X32 FILLCELL_253_544 ();
 FILLCELL_X32 FILLCELL_253_576 ();
 FILLCELL_X32 FILLCELL_253_608 ();
 FILLCELL_X32 FILLCELL_253_640 ();
 FILLCELL_X32 FILLCELL_253_672 ();
 FILLCELL_X32 FILLCELL_253_704 ();
 FILLCELL_X32 FILLCELL_253_736 ();
 FILLCELL_X32 FILLCELL_253_768 ();
 FILLCELL_X32 FILLCELL_253_800 ();
 FILLCELL_X32 FILLCELL_253_832 ();
 FILLCELL_X32 FILLCELL_253_864 ();
 FILLCELL_X32 FILLCELL_253_896 ();
 FILLCELL_X32 FILLCELL_253_928 ();
 FILLCELL_X32 FILLCELL_253_960 ();
 FILLCELL_X32 FILLCELL_253_992 ();
 FILLCELL_X32 FILLCELL_253_1024 ();
 FILLCELL_X32 FILLCELL_253_1056 ();
 FILLCELL_X32 FILLCELL_253_1088 ();
 FILLCELL_X32 FILLCELL_253_1120 ();
 FILLCELL_X32 FILLCELL_253_1152 ();
 FILLCELL_X32 FILLCELL_253_1184 ();
 FILLCELL_X32 FILLCELL_253_1216 ();
 FILLCELL_X32 FILLCELL_253_1248 ();
 FILLCELL_X32 FILLCELL_253_1280 ();
 FILLCELL_X32 FILLCELL_253_1312 ();
 FILLCELL_X32 FILLCELL_253_1344 ();
 FILLCELL_X32 FILLCELL_253_1376 ();
 FILLCELL_X32 FILLCELL_253_1408 ();
 FILLCELL_X32 FILLCELL_253_1440 ();
 FILLCELL_X32 FILLCELL_253_1472 ();
 FILLCELL_X32 FILLCELL_253_1504 ();
 FILLCELL_X32 FILLCELL_253_1536 ();
 FILLCELL_X32 FILLCELL_253_1568 ();
 FILLCELL_X32 FILLCELL_253_1600 ();
 FILLCELL_X32 FILLCELL_253_1632 ();
 FILLCELL_X32 FILLCELL_253_1664 ();
 FILLCELL_X32 FILLCELL_253_1696 ();
 FILLCELL_X32 FILLCELL_253_1728 ();
 FILLCELL_X32 FILLCELL_253_1760 ();
 FILLCELL_X32 FILLCELL_253_1792 ();
 FILLCELL_X32 FILLCELL_253_1824 ();
 FILLCELL_X32 FILLCELL_253_1856 ();
 FILLCELL_X8 FILLCELL_253_1888 ();
 FILLCELL_X1 FILLCELL_253_1896 ();
 FILLCELL_X32 FILLCELL_254_0 ();
 FILLCELL_X32 FILLCELL_254_32 ();
 FILLCELL_X32 FILLCELL_254_64 ();
 FILLCELL_X32 FILLCELL_254_96 ();
 FILLCELL_X32 FILLCELL_254_128 ();
 FILLCELL_X32 FILLCELL_254_160 ();
 FILLCELL_X32 FILLCELL_254_192 ();
 FILLCELL_X32 FILLCELL_254_224 ();
 FILLCELL_X32 FILLCELL_254_256 ();
 FILLCELL_X32 FILLCELL_254_288 ();
 FILLCELL_X32 FILLCELL_254_320 ();
 FILLCELL_X32 FILLCELL_254_352 ();
 FILLCELL_X32 FILLCELL_254_384 ();
 FILLCELL_X32 FILLCELL_254_416 ();
 FILLCELL_X32 FILLCELL_254_448 ();
 FILLCELL_X32 FILLCELL_254_480 ();
 FILLCELL_X32 FILLCELL_254_512 ();
 FILLCELL_X32 FILLCELL_254_544 ();
 FILLCELL_X32 FILLCELL_254_576 ();
 FILLCELL_X32 FILLCELL_254_608 ();
 FILLCELL_X32 FILLCELL_254_640 ();
 FILLCELL_X32 FILLCELL_254_672 ();
 FILLCELL_X32 FILLCELL_254_704 ();
 FILLCELL_X32 FILLCELL_254_736 ();
 FILLCELL_X32 FILLCELL_254_768 ();
 FILLCELL_X32 FILLCELL_254_800 ();
 FILLCELL_X32 FILLCELL_254_832 ();
 FILLCELL_X32 FILLCELL_254_864 ();
 FILLCELL_X32 FILLCELL_254_896 ();
 FILLCELL_X32 FILLCELL_254_928 ();
 FILLCELL_X32 FILLCELL_254_960 ();
 FILLCELL_X32 FILLCELL_254_992 ();
 FILLCELL_X32 FILLCELL_254_1024 ();
 FILLCELL_X32 FILLCELL_254_1056 ();
 FILLCELL_X32 FILLCELL_254_1088 ();
 FILLCELL_X32 FILLCELL_254_1120 ();
 FILLCELL_X32 FILLCELL_254_1152 ();
 FILLCELL_X32 FILLCELL_254_1184 ();
 FILLCELL_X32 FILLCELL_254_1216 ();
 FILLCELL_X32 FILLCELL_254_1248 ();
 FILLCELL_X32 FILLCELL_254_1280 ();
 FILLCELL_X32 FILLCELL_254_1312 ();
 FILLCELL_X32 FILLCELL_254_1344 ();
 FILLCELL_X32 FILLCELL_254_1376 ();
 FILLCELL_X32 FILLCELL_254_1408 ();
 FILLCELL_X32 FILLCELL_254_1440 ();
 FILLCELL_X32 FILLCELL_254_1472 ();
 FILLCELL_X32 FILLCELL_254_1504 ();
 FILLCELL_X32 FILLCELL_254_1536 ();
 FILLCELL_X32 FILLCELL_254_1568 ();
 FILLCELL_X32 FILLCELL_254_1600 ();
 FILLCELL_X32 FILLCELL_254_1632 ();
 FILLCELL_X32 FILLCELL_254_1664 ();
 FILLCELL_X32 FILLCELL_254_1696 ();
 FILLCELL_X32 FILLCELL_254_1728 ();
 FILLCELL_X32 FILLCELL_254_1760 ();
 FILLCELL_X32 FILLCELL_254_1792 ();
 FILLCELL_X32 FILLCELL_254_1824 ();
 FILLCELL_X32 FILLCELL_254_1856 ();
 FILLCELL_X8 FILLCELL_254_1888 ();
 FILLCELL_X1 FILLCELL_254_1896 ();
 FILLCELL_X32 FILLCELL_255_0 ();
 FILLCELL_X32 FILLCELL_255_32 ();
 FILLCELL_X32 FILLCELL_255_64 ();
 FILLCELL_X32 FILLCELL_255_96 ();
 FILLCELL_X32 FILLCELL_255_128 ();
 FILLCELL_X32 FILLCELL_255_160 ();
 FILLCELL_X32 FILLCELL_255_192 ();
 FILLCELL_X32 FILLCELL_255_224 ();
 FILLCELL_X32 FILLCELL_255_256 ();
 FILLCELL_X32 FILLCELL_255_288 ();
 FILLCELL_X32 FILLCELL_255_320 ();
 FILLCELL_X32 FILLCELL_255_352 ();
 FILLCELL_X32 FILLCELL_255_384 ();
 FILLCELL_X32 FILLCELL_255_416 ();
 FILLCELL_X32 FILLCELL_255_448 ();
 FILLCELL_X32 FILLCELL_255_480 ();
 FILLCELL_X32 FILLCELL_255_512 ();
 FILLCELL_X32 FILLCELL_255_544 ();
 FILLCELL_X32 FILLCELL_255_576 ();
 FILLCELL_X32 FILLCELL_255_608 ();
 FILLCELL_X32 FILLCELL_255_640 ();
 FILLCELL_X32 FILLCELL_255_672 ();
 FILLCELL_X32 FILLCELL_255_704 ();
 FILLCELL_X32 FILLCELL_255_736 ();
 FILLCELL_X32 FILLCELL_255_768 ();
 FILLCELL_X32 FILLCELL_255_800 ();
 FILLCELL_X32 FILLCELL_255_832 ();
 FILLCELL_X32 FILLCELL_255_864 ();
 FILLCELL_X32 FILLCELL_255_896 ();
 FILLCELL_X32 FILLCELL_255_928 ();
 FILLCELL_X32 FILLCELL_255_960 ();
 FILLCELL_X32 FILLCELL_255_992 ();
 FILLCELL_X32 FILLCELL_255_1024 ();
 FILLCELL_X32 FILLCELL_255_1056 ();
 FILLCELL_X32 FILLCELL_255_1088 ();
 FILLCELL_X32 FILLCELL_255_1120 ();
 FILLCELL_X32 FILLCELL_255_1152 ();
 FILLCELL_X32 FILLCELL_255_1184 ();
 FILLCELL_X32 FILLCELL_255_1216 ();
 FILLCELL_X32 FILLCELL_255_1248 ();
 FILLCELL_X32 FILLCELL_255_1280 ();
 FILLCELL_X32 FILLCELL_255_1312 ();
 FILLCELL_X32 FILLCELL_255_1344 ();
 FILLCELL_X32 FILLCELL_255_1376 ();
 FILLCELL_X32 FILLCELL_255_1408 ();
 FILLCELL_X32 FILLCELL_255_1440 ();
 FILLCELL_X32 FILLCELL_255_1472 ();
 FILLCELL_X32 FILLCELL_255_1504 ();
 FILLCELL_X32 FILLCELL_255_1536 ();
 FILLCELL_X32 FILLCELL_255_1568 ();
 FILLCELL_X32 FILLCELL_255_1600 ();
 FILLCELL_X32 FILLCELL_255_1632 ();
 FILLCELL_X32 FILLCELL_255_1664 ();
 FILLCELL_X32 FILLCELL_255_1696 ();
 FILLCELL_X32 FILLCELL_255_1728 ();
 FILLCELL_X32 FILLCELL_255_1760 ();
 FILLCELL_X32 FILLCELL_255_1792 ();
 FILLCELL_X32 FILLCELL_255_1824 ();
 FILLCELL_X32 FILLCELL_255_1856 ();
 FILLCELL_X8 FILLCELL_255_1888 ();
 FILLCELL_X1 FILLCELL_255_1896 ();
endmodule
